* SPICE NETLIST
***************************************

.SUBCKT TG A GND VDD G G_ Z
** N=6 EP=6 IP=0 FDC=2
M0 Z G A GND NM L=1.8e-07 W=2.2e-07 $X=-4200 $Y=-1655 $D=0
M1 Z G_ A VDD PM L=1.8e-07 W=2.2e-07 $X=-4200 $Y=500 $D=4
.ENDS
***************************************
