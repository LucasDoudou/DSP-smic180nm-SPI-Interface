* SPICE NETLIST
***************************************

.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=48
X0 1 2 3 4 10 11 9 Full_Adder_Sum $T=0 0 0 0 $X=10440 $Y=-19565
X1 5 6 7 8 10 11 12 Full_Adder_Sum $T=0 7690 0 0 $X=10440 $Y=-11875
.ENDS
***************************************
.SUBCKT 11FA B<0> B<1> B<2> B<3> B<4> B<5> A<0> A<1> A<2> A<3> A<4> A<5> S<1> S<2> S<3> S<4> S<5> S<0> B<9> A<7>
+ A<8> B<10> A<6> B<6> A<9> A<10> B<8> B<7> S<6> S<7> S<8> S<9> S<10> COUT GND VDD
** N=68 EP=36 IP=133 FDC=308
X0 58 GND VDD S<0> 38 45 ICV_1 $T=31380 -61685 0 0 $X=27265 $Y=-58600
X1 59 GND VDD S<1> 39 46 ICV_1 $T=31380 -53995 0 0 $X=27265 $Y=-50910
X2 60 GND VDD S<2> 40 47 ICV_1 $T=31380 -46120 0 0 $X=27265 $Y=-43035
X3 61 GND VDD S<3> 41 44 ICV_1 $T=31380 -38430 0 0 $X=27265 $Y=-35345
X4 62 GND VDD S<4> 42 48 ICV_1 $T=31380 -30605 0 0 $X=27265 $Y=-27520
X5 63 GND VDD S<5> 43 37 ICV_1 $T=31380 -22915 0 0 $X=27265 $Y=-19830
X6 64 GND VDD S<6> 49 54 ICV_1 $T=51680 -53805 0 0 $X=47565 $Y=-50720
X7 65 GND VDD S<7> 50 55 ICV_1 $T=51680 -46115 0 0 $X=47565 $Y=-43030
X8 66 GND VDD S<8> 51 56 ICV_1 $T=51680 -38240 0 0 $X=47565 $Y=-35155
X9 67 GND VDD S<9> 52 57 ICV_1 $T=51680 -30550 0 0 $X=47565 $Y=-27465
X10 68 GND VDD S<10> 53 COUT ICV_1 $T=51680 -22915 0 0 $X=47565 $Y=-19830
X11 57 A<10> B<10> 53 GND VDD 68 Full_Adder_Sum $T=22055 -265 0 0 $X=32495 $Y=-19830
X12 GND A<0> B<0> 38 45 A<1> B<1> 39 58 GND VDD 59 ICV_2 $T=1755 -39035 0 0 $X=12195 $Y=-58600
X13 46 A<2> B<2> 40 47 A<3> B<3> 41 60 GND VDD 61 ICV_2 $T=1755 -23470 0 0 $X=12195 $Y=-43035
X14 44 A<4> B<4> 42 48 A<5> B<5> 43 62 GND VDD 63 ICV_2 $T=1755 -7955 0 0 $X=12195 $Y=-27520
X15 37 A<6> B<6> 49 54 A<7> B<7> 50 64 GND VDD 65 ICV_2 $T=22055 -31155 0 0 $X=32495 $Y=-50720
X16 55 A<8> B<8> 51 56 A<9> B<9> 52 66 GND VDD 67 ICV_2 $T=22055 -15590 0 0 $X=32495 $Y=-35155
.ENDS
***************************************
.SUBCKT And_Gate VIN_B VIN_A VDD GND VOUT
** N=7 EP=5 IP=0 FDC=6
M0 6 VIN_A 7 GND NM L=1.8e-07 W=2.2e-07 $X=1890 $Y=-4485 $D=0
M1 GND VIN_B 6 GND NM L=1.8e-07 W=2.2e-07 $X=2690 $Y=-4485 $D=0
M2 VOUT 7 GND GND NM L=1.8e-07 W=2.2e-07 $X=3490 $Y=-4485 $D=0
M3 7 VIN_A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1890 $Y=-2095 $D=4
M4 VDD VIN_B 7 VDD PM L=1.8e-07 W=4.4e-07 $X=2610 $Y=-2095 $D=4
M5 VOUT 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3330 $Y=-2095 $D=4
.ENDS
***************************************
.SUBCKT 6_AND_test Y<0> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND Z<0> A<0> A<1> A<2> A<3> A<4>
** N=15 EP=15 IP=30 FDC=36
X0 X<0> Y<0> VDD GND Z<0> And_Gate $T=2375 -2105 0 0 $X=3355 $Y=-7730
X1 X<1> Y<0> VDD GND A<0> And_Gate $T=5555 -2105 0 0 $X=6535 $Y=-7730
X2 X<2> Y<0> VDD GND A<1> And_Gate $T=8735 -2105 0 0 $X=9715 $Y=-7730
X3 X<3> Y<0> VDD GND A<2> And_Gate $T=11915 -2105 0 0 $X=12895 $Y=-7730
X4 X<4> Y<0> VDD GND A<3> And_Gate $T=15095 -2105 0 0 $X=16075 $Y=-7730
X5 X<5> Y<0> VDD GND A<4> And_Gate $T=18275 -2105 0 0 $X=19255 $Y=-7730
.ENDS
***************************************
.SUBCKT 6_FA_v3 S<0> S<1> S<2> S<3> S<4> S<5> S<6> GND A<0> B<0> A<1> B<1> A<2> B<2> A<3> B<3> A<4> B<4> A<5> B<5>
+ VDD
** N=38 EP=21 IP=78 FDC=168
X0 33 GND VDD S<0> 22 29 ICV_1 $T=11635 -18360 0 0 $X=7520 $Y=-15275
X1 34 GND VDD S<1> 23 30 ICV_1 $T=11635 -10670 0 0 $X=7520 $Y=-7585
X2 35 GND VDD S<2> 24 31 ICV_1 $T=11635 -2795 0 0 $X=7520 $Y=290
X3 36 GND VDD S<3> 25 28 ICV_1 $T=11635 4895 0 0 $X=7520 $Y=7980
X4 37 GND VDD S<4> 26 32 ICV_1 $T=11635 12720 0 0 $X=7520 $Y=15805
X5 38 GND VDD S<5> 27 S<6> ICV_1 $T=11635 20410 0 0 $X=7520 $Y=23495
X6 GND A<0> B<0> 22 GND VDD 33 Full_Adder_Sum $T=-17990 4290 0 0 $X=-7550 $Y=-15275
X7 29 A<1> B<1> 23 GND VDD 34 Full_Adder_Sum $T=-17990 11980 0 0 $X=-7550 $Y=-7585
X8 30 A<2> B<2> 24 GND VDD 35 Full_Adder_Sum $T=-17990 19855 0 0 $X=-7550 $Y=290
X9 31 A<3> B<3> 25 GND VDD 36 Full_Adder_Sum $T=-17990 27545 0 0 $X=-7550 $Y=7980
X10 28 A<4> B<4> 26 GND VDD 37 Full_Adder_Sum $T=-17990 35370 0 0 $X=-7550 $Y=15805
X11 32 A<5> B<5> 27 GND VDD 38 Full_Adder_Sum $T=-17990 43060 0 0 $X=-7550 $Y=23495
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=12
X0 1 3 4 5 6 And_Gate $T=0 0 0 0 $X=980 $Y=-5625
X1 2 3 4 5 7 And_Gate $T=3180 0 0 0 $X=4160 $Y=-5625
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=24
X0 1 2 7 6 5 8 9 ICV_3 $T=0 0 0 0 $X=980 $Y=-5625
X1 3 4 10 6 5 11 12 ICV_3 $T=6360 0 0 0 $X=7340 $Y=-5625
.ENDS
***************************************
.SUBCKT 5_6_Multiplier X<0> X<1> X<2> X<3> X<4> X<5> Y<1> Y<0> Z<0> Z<1> GND Y<3> Y<4> Y<2> Z<2> Z<3> Z<4> Z<5> Z<6> Z<7>
+ Z<8> Z<9> Z<10> VDD
** N=88 EP=24 IP=222 FDC=852
X0 83 GND VDD Z<1> 54 61 ICV_1 $T=48685 -77935 0 0 $X=44570 $Y=-74850
X1 84 GND VDD 33 55 62 ICV_1 $T=48685 -70245 0 0 $X=44570 $Y=-67160
X2 85 GND VDD 34 56 63 ICV_1 $T=48685 -62370 0 0 $X=44570 $Y=-59285
X3 86 GND VDD 36 57 60 ICV_1 $T=48685 -54680 0 0 $X=44570 $Y=-51595
X4 87 GND VDD 32 58 64 ICV_1 $T=48685 -46855 0 0 $X=44570 $Y=-43770
X5 88 GND VDD 35 59 31 ICV_1 $T=48685 -39165 0 0 $X=44570 $Y=-36080
X6 GND 49 25 54 GND VDD 83 Full_Adder_Sum $T=19060 -55285 0 0 $X=29500 $Y=-74850
X7 61 50 26 55 GND VDD 84 Full_Adder_Sum $T=19060 -47595 0 0 $X=29500 $Y=-67160
X8 62 51 27 56 GND VDD 85 Full_Adder_Sum $T=19060 -39720 0 0 $X=29500 $Y=-59285
X9 63 52 28 57 GND VDD 86 Full_Adder_Sum $T=19060 -32030 0 0 $X=29500 $Y=-51595
X10 60 53 29 58 GND VDD 87 Full_Adder_Sum $T=19060 -24205 0 0 $X=29500 $Y=-43770
X11 64 GND 30 59 GND VDD 88 Full_Adder_Sum $T=19060 -16515 0 0 $X=29500 $Y=-36080
X12 Y<2> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 65 66 67 68 69 70 6_AND_test $T=51110 -22420 0 0 $X=54270 $Y=-30150
X13 Y<3> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 71 72 73 74 75 76 6_AND_test $T=75810 -22420 0 0 $X=78970 $Y=-30150
X14 Y<4> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 77 78 79 80 81 82 6_AND_test $T=100535 -22420 0 0 $X=103695 $Y=-30150
X15 Z<2> 41 40 38 39 42 37 GND 33 65 34 66 36 67 32 68 35 69 31 70
+ VDD
+ 6_FA_v3 $T=62150 -60875 0 0 $X=53915 $Y=-76150
X16 Z<3> 44 46 45 47 48 43 GND 41 71 40 72 38 73 39 74 42 75 37 76
+ VDD
+ 6_FA_v3 $T=86850 -60875 0 0 $X=78615 $Y=-76150
X17 Z<4> Z<5> Z<6> Z<7> Z<8> Z<9> Z<10> GND 44 77 46 78 45 79 47 80 48 81 43 82
+ VDD
+ 6_FA_v3 $T=111575 -60875 0 0 $X=103340 $Y=-76150
X18 X<0> X<1> X<2> X<3> GND VDD Y<1> 25 26 Y<1> 27 28 ICV_4 $T=18540 -72855 0 90 $X=19065 $Y=-71875
X19 X<4> X<5> X<0> X<1> GND VDD Y<1> 29 30 Y<0> Z<0> 49 ICV_4 $T=18540 -60135 0 90 $X=19065 $Y=-59155
X20 X<2> X<3> X<4> X<5> GND VDD Y<0> 50 51 Y<0> 52 53 ICV_4 $T=18540 -47415 0 90 $X=19065 $Y=-46435
.ENDS
***************************************
.SUBCKT DSP_final_v1 C<0> C<4> C<3> C<2> C<5> C<1> C<8> C<6> C<7> C<10> C<9> A<2> A<0> A<4> A<1> A<3> A<5> GND D<0> B<0>
+ D<1> B<1> D<2> B<2> D<3> B<3> VDD P<0> P<4> P<3> P<2> P<5> P<1> P<10> P<9> P<11> P<6> P<7> P<8>
** N=66 EP=39 IP=120 FDC=1272
X0 31 GND VDD 32 inv $T=141520 -3830 0 270 $X=144605 $Y=-1715
X1 51 GND VDD 30 inv $T=141520 -2330 0 270 $X=144605 $Y=-215
X2 33 GND VDD 35 inv $T=149210 -3830 0 270 $X=152295 $Y=-1715
X3 52 GND VDD 29 inv $T=149210 -2330 0 270 $X=152295 $Y=-215
X4 36 GND VDD 39 inv $T=157085 -3830 0 270 $X=160170 $Y=-1715
X5 53 GND VDD 34 inv $T=157085 -2330 0 270 $X=160170 $Y=-215
X6 40 GND VDD 38 inv $T=164775 -3830 0 270 $X=167860 $Y=-1715
X7 54 GND VDD 37 inv $T=164775 -2330 0 270 $X=167860 $Y=-215
X8 GND D<0> B<0> 31 GND VDD 51 Full_Adder_Sum $T=164170 27295 0 270 $X=144605 $Y=3040
X9 32 D<1> B<1> 33 GND VDD 52 Full_Adder_Sum $T=171860 27295 0 270 $X=152295 $Y=3040
X10 35 D<2> B<2> 36 GND VDD 53 Full_Adder_Sum $T=179735 27295 0 270 $X=160170 $Y=3040
X11 39 D<3> B<3> 40 GND VDD 54 Full_Adder_Sum $T=187425 27295 0 270 $X=167860 $Y=3040
X12 C<0> C<1> C<2> C<3> C<4> C<5> 3 1 5 4 6 7 P<1> P<2> P<3> P<4> P<5> P<0> C<9> 8
+ 9 C<10> 2 C<6> 11 10 C<8> C<7> P<6> P<7> P<8> P<9> P<10> P<11> GND VDD
+ 11FA $T=54410 44955 1 270 $X=67075 $Y=-6830
X13 A<0> A<1> A<2> A<3> A<4> A<5> 29 30 3 1 GND 37 38 34 5 4 6 7 2 8
+ 9 11 10 VDD
+ 5_6_Multiplier $T=52050 20650 0 0 $X=67615 $Y=-55500
.ENDS
***************************************
