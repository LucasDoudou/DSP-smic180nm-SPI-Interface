//*Spectre Model Format
simulator lang=spectre  insensitive=yes
// *
// *
// * no part of this file can be released without the consent of smic.
// *
// *******************************************************************************************
// * 0.18um mixed signal 1p6m with mim salicide 1.8v/3.3v rf spice model (for spectre only)  *
// *******************************************************************************************
// *
// * release version    : 1.6
// *
// * release date       : 07/02/2007
// *
// * simulation tool    : Cadence spectre V6.0
// *
// * model type         :
// *   mosfet           : bsim3v3.2
// *   junction diode   : spectre level 1
// *
// * model and subcircuit name         :
// *   mosfet           :
//*        *------------------------------------------*
//*        |     MOSFET model   |   1.8V   |   3.3V   |
//*        |==========================================|
//*        |        NMOS        |  n18_rf  |  n33_rf  |
//*        *------------------------------------------*
//*        |       DNWMOS       | dnw18_rf | dnw33_rf |
//*        *------------------------------------------*
//*        |        PMOS        |  p18_rf  |  p33_rf  |
//*        *------------------------------------------*
//*
//*        *--------------------------------------------------*
//*        |     MOSFET subckt  |     1.8V     |    3.3V      |
//*        |==================================================|
//*        |        NMOS        |  n18_ckt_rf  |  n33_ckt_rf  |
//*        *--------------------------------------------------*
//*        |       DNWMOS       | dnw18_ckt_rf | dnw33_ckt_rf |
//*        *--------------------------------------------------*
//*        |        PMOS        |  p18_ckt_rf  |  p33_ckt_rf  |
//*        *--------------------------------------------------*
//*
//*************************
//* 1.8V RF NMOS Subcircuit
//*************************
//* 1=drain, 2=gate, 3=source, 4=bulk
//* lr=gate length, wr=finger width, nf=finger number
subckt n18_ckt_rf (1 2 3 4) 
//* scalable unit parameter
//* euqivalent circuit saclable parameter
parameters lr=0.18u wr=10u nf=2
+rdc_n18      = max(17*(1/(pow(wr*1e6,0.9))), 1e-3)
+rsc_n18      = max(17*(1/(pow(wr*1e6,0.9))), 1e-3)
+cgdo_n18     = max((0+dcgdo_n18_rf), 0)
+cgso_n18     = max((0+dcgso_n18_rf), 0)
//*****************************************
lgate       (2 20)  inductor   l=1p
rgate       (20 21) resistor   r=max((1542.7*lr*1e6+165.64)*pow(wr*1e6,-0.9019*lr*1e6-0.5975)*pow(nf,-0.9912*pow(wr*1e6,-0.1348)), 1e-3)
cgd_ext     (20 11) capacitor  c=max(((8.85e-16*lr*lr*1e12-4.83e-16*lr*1e6+3.92e-16)*wr*1e6+2.95e-16)*nf+3.19e-16*pow(wr*1e6,0.402), 1e-18)
cgs_ext     (20 31) capacitor  c=max(((4.82e-16*lr*1e6+9.58e-17)*pow(wr*1e6,2.3513*lr*1e6-1.3178))*nf+1.34e-15*pow(wr*1e6,-0.763), 1e-18)
cds_ext     (15 31) capacitor  c=max(((3.37e-17*pow(lr*1e6,-1.38))*wr*1e6+1.89e-16)*nf+(-1.21e-14*lr*lr*1e12+9.83e-15*lr*1e6-9.86e-16)*pow(wr*1e6,0.505), 1e-18)
rds         (11 15) resistor   r=0.01
ldrain      (1 11)  inductor   l=1p
lsource     (3 31)  inductor   l=1p
//*****************************************
djdb (12 11) ndio18_rf area=(nf/2*(0.8-2*0.07)*wr*1e6)*1e-12 pj=(-0.048*log(wr*1e6)+1.1121)*(nf*wr)
djsb (32 31) ndio18_rf area=((nf/2-1)*(0.8-2*0.07)*wr*1e6+(0.8-0.07)*wr*1e6*2)*1e-12 pj=(-0.0567*log(wr*1e6)+1.1608)*(nf*wr)
//*****************************************
rsub1      (41  4)  resistor   r=max(341.64*pow(nf,-0.5321), 1e-3)
rsub2      (41  12) resistor   r=max(341.64*pow(nf,-0.5321), 1e-3)
rsub3      (41  32) resistor   r=12000
//* --------- ideal mos transistor ----------------------
main (11 21 31 41) n18_rf l=lr w=wr m=nf ad = 0 as = 0 pd = 0 ps = 0
// * mos model
model n18_rf bsim3v3 {
1: type=n
// * general parameters
// *
+lmin = 1.6e-7 lmax = 5.2e-7 wmin = 4.8e-7 
+wmax = 1.002e-5 tnom = 25.0 version = 3.2 
+tox = 3.87e-09+dtox_n18_rf toxm = 3.87e-09 xj = 1.6000000e-07 
+nch = 3.8694000e+17 lln = 1.1205959 lwn = 0.9200000 
+wln = 1.0599999 wwn = 0.8768474 lint = 1.5757085e-08 
+ll = 2.6352781e-16 lw = -2.2625584e-16 lwl = -2.0576711e-22 
+wint = -1.4450482e-09 wl = -2.3664573e-16 ww = -3.6409690e-14 
+wwl = -4.0000000e-21 mobmod = 1 binunit = 2 
+xl = 1.8e-8+dxl_n18_rf xw = 0.00+dxw_n18_rf dwg = -5.9600000e-09 
+dwb = 4.5000000e-09 
// * diode parameters
+dskip = no ldif = 7.00e-08 hdif = 2.00e-07 
+rsh = 7.08 rd = 0 rs = 0 
+rsc = rsc_n18 rdc = rdc_n18 
// *
// * threshold voltage parameters
// *
+vth0 = 0.39+dvth_n18_rf wvth0 = -2.9709472e-08 pvth0 = 5.0000000e-16+dpvth0_n18_rf 
+k1 = 0.6801043 wk1 = -2.4896840e-08 pk1 = 1.3000000e-15 
+k2 = -4.9977830e-02 k3 = 10.0000000 dvt0 = 1.3000000 
+dvt1 = 0.5771635 dvt2 = -0.1717554 dvt0w = 0.00 
+dvt1w = 0.00 dvt2w = 0.00 nlx = 7.5451030e-08 
+w0 = 5.5820150e-07 k3b = -3.0000000 
// *
// * mobility parameters
// *
+vsat = 8.2500000e+04 pvsat = -8.3000000e-10 ua = -1.0300000e-09 
+lua = 7.7349790e-19 pua = -1.0000000e-24 ub = 2.3666682e-18 
+uc = 1.2000000e-10 puc = 1.5000000e-24 rdsw = 55.5497200 
+prwb = -0.2400000 prwg = 0.4000000 wr = 1.0000000 
+u0 = 3.4000000e-02 lu0 = 2.3057663e-11 wu0 = -3.1009695e-09 
+a0 = 0.8300000 keta = -3.0000000e-03 lketa = -1.7000000e-09 
+a1 = 0.00 a2 = 0.9900000 ags = 0.3200000 
+b0 = 6.0000000e-08 b1 = 0.00 
// *
// * subthreshold current parameters
// *
+voff = -0.1030000 lvoff = -3.3000000e-09 nfactor = 1.2500000 
+lnfactor = 4.5000000e-08 cit = 0.00 cdsc = 0.00 
+cdscb = 0.00 cdscd = 1.0000000e-04 eta0 = 2.8000001e-02 
+etab = -2.7000001e-02 dsub = 0.4000000 
// *
// * rout parameters
// *
+pclm = 1.2000000 ppclm = 2.9999999e-15 pdiblc1 = 2.5000000e-02 
+pdiblc2 = 3.8000000e-03 ppdiblc2 = 2.7000001e-16 pdiblcb = 0.00 
+drout = 0.5600000 pscbe1 = 3.4500000e+08 pscbe2 = 1.0000000e-06 
+pvag = 0.00 delta = 1.0000000e-02 alpha0 = 1.7753978e-08 
+alpha1 = 0.1764000 lalpha1 = 7.6250000e-09 beta0 = 11.1683940 
// *
// * temperature effects parameters
// *
+kt1 = -0.2572866 kt2 = -4.0000000e-02 at = 3.7000000e+04 
+pat = -7.5000000e-10 ute = -1.5500000 ua1 = 1.7600000e-09 
+lua1 = 6.0000000e-18 wua1 = -1.1000000e-16 pua1 = -5.0000000e-25 
+ub1 = -2.4000000e-18 uc1 = -1.0000000e-10 luc1 = 1.6999999e-17 
+puc1 = -3.0000000e-24 kt1l = -1.0000000e-09 prt = -55.0000000 
// *
// * capacitance parameters
// *
+cj = 0 mj = 0.346 pb = 0.7 
+cjsw = 0 mjsw = 0.538 pbsw = 1 
+cjswg = 0 mjswg = 0.538 pbswg = 1 
+tcj = 8.42e-04 tcjsw = 6.69e-04 tcjswg = 6.69e-04 
+tpb = 1.47e-03 tpbsw = 8.68e-04 tpbswg = 8.68e-04 
+js = 3.52e-07 jsw = 3.0e-13 n = 1.0392 
+xti = 3.25 nqsmod = 0 elm = 5 
+cgdo = cgdo_n18 cgso = cgso_n18 tlevc = 1 
+capmod = 3 xpart = 1 cf = 0.00 
+acde = 0.64 moin = 24 noff = 1.2025 
+dlc = 8.5e-09 dwc = 4.5e-08 
+noimod  = 1 flkmod = 1 af = 0.85 kf = 1.5e-24 
}
// * junction diode model
model ndio18_rf diode
+is = 3.52e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15 
+n = 1.0233 ns = 1.0233  ik = 1.52e+05 ikp = 4.32e-04 
+bv = 11.0 ibv = 277.78 
+trs = 1.51e-03 eg = 1.16 tnom = 25.0  xti = 3.0
+rs = 8.89e-09 
+cjo = 9.68e-04+dcj_n18_rf
+cjsw = 4.18e-10+dcjsw_n18_rf 
+mj = 0.346 vj = 0.7  mjsw = 0.538 
+vjsw = 1 cta = 0.000842 ctp = 0.000669 
+pta = 0.00147 ptp = 0.000868 tlev = 1 
+tlevc = 1 fc = 0 
ends n18_ckt_rf
//***************************
//* 1.8V RF DNWMOS Subcircuit
//***************************
//* 1=drain, 2=gate, 3=source, 4=bulk, 5=DNW
//* lr=gate length, wr=finger width, nf=finger number, laddr=DNW diode add length, waddr=DNW didoe add width
subckt dnw18_ckt_rf (1 2 3 4 5) 
//* scalable unit parameter
//* euqivalent circuit saclable parameter
parameters lr=0.18u wr=10u nf=2 laddr=10u waddr=10u
+rdc_n18      = max(17*(1/(pow(wr*1e6,0.9))), 1e-3)
+rsc_n18      = max(17*(1/(pow(wr*1e6,0.9))), 1e-3)
+cgdo_n18     = max((0+dcgdo_n18_rf), 0)
+cgso_n18     = max((0+dcgso_n18_rf), 0)
//*****************************************
lgate       (2 20)  inductor   l=1p
rgate       (20 21) resistor   r=max((1542.7*lr*1e6+165.64)*pow(wr*1e6,-0.9019*lr*1e6-0.5975)*pow(nf,-0.9912*pow(wr*1e6,-0.1348)), 1e-3)
cgd_ext     (20 11) capacitor  c=max(((8.85e-16*lr*lr*1e12-4.83e-16*lr*1e6+3.92e-16)*wr*1e6+2.95e-16)*nf+3.19e-16*pow(wr*1e6,0.402), 1e-18)
cgs_ext     (20 31) capacitor  c=max(((4.82e-16*lr*1e6+9.58e-17)*pow(wr*1e6,2.3513*lr*1e6-1.3178))*nf+1.34e-15*pow(wr*1e6,-0.763), 1e-18)
cds_ext     (15 31) capacitor  c=max(((3.37e-17*pow(lr*1e6,-1.38))*wr*1e6+1.89e-16)*nf+(-1.21e-14*lr*lr*1e12+9.83e-15*lr*1e6-9.86e-16)*pow(wr*1e6,0.505), 1e-18)
rds         (11 15) resistor   r=0.01
ldrain      (1 11)  inductor   l=1p
lsource     (3 31)  inductor   l=1p
//*****************************************
djdb (12 11) ndio18_rf area=(nf/2*(0.8-2*0.07)*wr*1e6)*1e-12 pj=(-0.048*log(wr*1e6)+1.1121)*(nf*wr)
djsb (32 31) ndio18_rf area=((nf/2-1)*(0.8-2*0.07)*wr*1e6+(0.8-0.07)*wr*1e6*2)*1e-12 pj=(-0.0567*log(wr*1e6)+1.1608)*(nf*wr)
djdnw (4 5) diobpw_rf area=(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+2*laddr)*(wr+2*waddr) pj=2*(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+wr+2*(laddr+waddr))
//*****************************************
rsub1      (41  4)  resistor   r=max(341.64*pow(nf,-0.5321), 1e-3)
rsub2      (41  12) resistor   r=max(341.64*pow(nf,-0.5321), 1e-3)
rsub3      (41  32) resistor   r=12000
//* --------- ideal mos transistor ----------------------
main (11 21 31 41) dnw18_rf l=lr w=wr m=nf ad = 0 as = 0 pd = 0 ps = 0
// * mos model
model dnw18_rf bsim3v3 {
1: type=n
// * general parameters
// *
+lmin = 1.6e-7 lmax = 5.2e-7 wmin = 4.8e-7 
+wmax = 1.002e-5 tnom = 25.0 version = 3.2 
+tox = 3.87e-09+dtox_n18_rf toxm = 3.87e-09 xj = 1.6000000e-07 
+nch = 3.8694000e+17 lln = 1.1205959 lwn = 0.9200000 
+wln = 1.0599999 wwn = 0.8768474 lint = 1.5757085e-08 
+ll = 2.6352781e-16 lw = -2.2625584e-16 lwl = -2.0576711e-22 
+wint = -1.4450482e-09 wl = -2.3664573e-16 ww = -3.6409690e-14 
+wwl = -4.0000000e-21 mobmod = 1 binunit = 2 
+xl = 1.8e-8+dxl_n18_rf xw = 0.00+dxw_n18_rf dwg = -5.9600000e-09 
+dwb = 4.5000000e-09 
// * diode parameters
+dskip = no ldif = 7.00e-08 hdif = 2.00e-07 
+rsh = 7.08 rd = 0 rs = 0 
+rsc = rsc_n18 rdc = rdc_n18 
// *
// * threshold voltage parameters
// *
+vth0 = 0.39+dvth_n18_rf wvth0 = -2.9709472e-08 pvth0 = 5.0000000e-16+dpvth0_n18_rf 
+k1 = 0.6801043 wk1 = -2.4896840e-08 pk1 = 1.3000000e-15 
+k2 = -4.9977830e-02 k3 = 10.0000000 dvt0 = 1.3000000 
+dvt1 = 0.5771635 dvt2 = -0.1717554 dvt0w = 0.00 
+dvt1w = 0.00 dvt2w = 0.00 nlx = 7.5451030e-08 
+w0 = 5.5820150e-07 k3b = -3.0000000 
// *
// * mobility parameters
// *
+vsat = 8.2500000e+04 pvsat = -8.3000000e-10 ua = -1.0300000e-09 
+lua = 7.7349790e-19 pua = -1.0000000e-24 ub = 2.3666682e-18 
+uc = 1.2000000e-10 puc = 1.5000000e-24 rdsw = 55.5497200 
+prwb = -0.2400000 prwg = 0.4000000 wr = 1.0000000 
+u0 = 3.4000000e-02 lu0 = 2.3057663e-11 wu0 = -3.1009695e-09 
+a0 = 0.8300000 keta = -3.0000000e-03 lketa = -1.7000000e-09 
+a1 = 0.00 a2 = 0.9900000 ags = 0.3200000 
+b0 = 6.0000000e-08 b1 = 0.00 
// *
// * subthreshold current parameters
// *
+voff = -0.1030000 lvoff = -3.3000000e-09 nfactor = 1.2500000 
+lnfactor = 4.5000000e-08 cit = 0.00 cdsc = 0.00 
+cdscb = 0.00 cdscd = 1.0000000e-04 eta0 = 2.8000001e-02 
+etab = -2.7000001e-02 dsub = 0.4000000 
// *
// * rout parameters
// *
+pclm = 1.2000000 ppclm = 2.9999999e-15 pdiblc1 = 2.5000000e-02 
+pdiblc2 = 3.8000000e-03 ppdiblc2 = 2.7000001e-16 pdiblcb = 0.00 
+drout = 0.5600000 pscbe1 = 3.4500000e+08 pscbe2 = 1.0000000e-06 
+pvag = 0.00 delta = 1.0000000e-02 alpha0 = 1.7753978e-08 
+alpha1 = 0.1764000 lalpha1 = 7.6250000e-09 beta0 = 11.1683940 
// *
// * temperature effects parameters
// *
+kt1 = -0.2572866 kt2 = -4.0000000e-02 at = 3.7000000e+04 
+pat = -7.5000000e-10 ute = -1.5500000 ua1 = 1.7600000e-09 
+lua1 = 6.0000000e-18 wua1 = -1.1000000e-16 pua1 = -5.0000000e-25 
+ub1 = -2.4000000e-18 uc1 = -1.0000000e-10 luc1 = 1.6999999e-17 
+puc1 = -3.0000000e-24 kt1l = -1.0000000e-09 prt = -55.0000000 
// *
// * capacitance parameters
// *
+cj = 0 mj = 0.346 pb = 0.7 
+cjsw = 0 mjsw = 0.538 pbsw = 1 
+cjswg = 0 mjswg = 0.538 pbswg = 1 
+tcj = 8.42e-04 tcjsw = 6.69e-04 tcjswg = 6.69e-04 
+tpb = 1.47e-03 tpbsw = 8.68e-04 tpbswg = 8.68e-04 
+js = 3.52e-07 jsw = 3.0e-13 n = 1.0392 
+xti = 3.25 nqsmod = 0 elm = 5 
+cgdo = cgdo_n18 cgso = cgso_n18 tlevc = 1 
+capmod = 3 xpart = 1 cf = 0.00 
+acde = 0.64 moin = 24 noff = 1.2025 
+dlc = 8.5e-09 dwc = 4.5e-08 
+noimod  = 1 flkmod = 1 af = 0.85 kf = 1.5e-24 
}
// * junction diode model
model ndio18_rf diode
+is = 3.52e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15 
+n = 1.0233 ns = 1.0233  ik = 1.52e+05 ikp = 4.32e-04 
+bv = 11.0 ibv = 277.78 
+trs = 1.51e-03 eg = 1.16 tnom = 25.0  xti = 3.0
+rs = 8.89e-09 
+cjo = 9.68e-04+dcj_n18_rf
+cjsw = 4.18e-10+dcjsw_n18_rf 
+mj = 0.346 vj = 0.7  mjsw = 0.538 
+vjsw = 1 cta = 0.000842 ctp = 0.000669 
+pta = 0.00147 ptp = 0.000868 tlev = 1 
+tlevc = 1 fc = 0 
// * DNW junction diode model
model diobpw_rf diode
+level = 1 is = 1.50e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1.00e-15 
+n = 1.0213 ns = 1.0213 rs = 2.51e-08 ik = 2.40e+05 ikp = 1.60E-03 
+bv = 15.0 ibv = 1.04e+02 
+trs = 1.77e-03 cta = 0.0012 ctp = 0.00107 
+eg = 1.16 tnom = 25.0 pta = 0.0019 
+ptp = 0.00193 xti = 3.0 cjo = 0.000536 
+mj = 0.343 vj = 0.693 cjsw = 3.22e-10 
+mjsw = 0.361 vjsw = 0.715 tlev = 1 
+tlevc = 1 area = 9.6e-9 perim = 4e-4 
+fc = 0 
ends dnw18_ckt_rf
//*************************
//* 1.8V RF PMOS Subcircuit
//*************************
//* 1=drain, 2=gate, 3=source, 4=bulk
//* lr=gate length, wr=finger width, nf=finger number
subckt p18_ckt_rf (1 2 3 4) 
//* scalable unit parameter
//* euqivalent circuit saclable parameter
parameters lr=0.18u wr=10u nf=2
+cgdo_p18     = max((0+dcgdo_p18_rf), 0)
+cgso_p18     = max((0+dcgso_p18_rf), 0)
//*****************************************
lgate       (2 20)  inductor   l=1p
rgate       (20 21) resistor   r=max((9852.3*lr*1e6-654.92)*pow(wr*1e6,7.3896*lr*lr*1e12-5.4762*lr*1e6-0.0697)*pow(nf,-1.0664*pow(wr*1e6,2.8625*lr*lr*1e12-1.919*lr*1e6+0.2309)), 1e-3)
cgd_ext     (20 11) capacitor  c=max(((4.03e-16*lr*1e6+3.02e-16)*wr*1e6+3.06e-16)*nf+2.94e-16*pow(wr*1e6,0.373), 1e-18)
cgs_ext     (20 31) capacitor  c=max((1.10e-15*pow(wr*1e6,-0.367))*nf+(-1.06e-15*log(wr*1e6)+2.55e-15), 1e-18)
cds_ext     (15 31) capacitor  c=max((3.46e-16*wr*1e6+2.44e-16)*nf+(6.79e-17*wr*wr*1e12-3.13e-16*wr*1e6+1.17e-15), 1e-18)
rds         (11 15) resistor   r=0.01
ldrain      (1 11)  inductor   l=1p
lsource     (3 31)  inductor   l=1p
//*****************************************
djdb (11 12) pdio18_rf area=(nf/2*(0.8-2*0.07)*wr*1e6)*1e-12 pj=(-0.0492*log(wr*1e6)+1.1146)*(nf*wr)
djsb (31 32) pdio18_rf area=((nf/2-1)*(0.8-2*0.07)*wr*1e6+(0.8-0.07)*wr*1e6*2)*1e-12 pj=(-0.0582*log(wr*1e6)+1.1649)*(nf*wr)
//*****************************************
rsub1      (41  4)  resistor   r=max(241.1*pow(nf,-0.4726), 1e-3)
rsub2      (41  12) resistor   r=max(241.1*pow(nf,-0.4726), 1e-3)
rsub3      (41  32) resistor   r=18000
//* --------- ideal mos transistor ----------------------
main (11 21 31 41) p18_rf l=lr w=wr m=nf ad = 0 as = 0 pd = 0 ps = 0
// * mos model
model p18_rf bsim3v3 {
1: type=p
// * general parameters
// *
+lmin = 1.6e-7 lmax = 5.2e-7 wmin = 4.8e-7 
+wmax = 1.002e-5 tnom = 25.0 version = 3.2 
+tox = 3.74e-09+dtox_p18_rf toxm = 3.74e-09 xj = 1.7000001e-07 
+nch = 5.5000000e+17 lln = 1.0000000 lwn = 1.0000000 
+wln = 1.0450000 wwn = 1.0000000 lint = 1.0000000e-08 
+ll = 3.4000000e-15 lw = -3.3600000e-16 lwl = 0.00 
+wint = 8.0000010e-09 wl = 3.5904200e-15 ww = -1.8999999e-15 
+wwl = -1.1205000e-21 mobmod = 1 binunit = 2 
+xl = -5.7e-09+dxl_p18_rf xw = 0.00+dxw_p18_rf dwg = -1.7361970e-08 
+dwb = 2.0000000e-08 
// * diode parameters
+dskip = no ldif = 7.00e-08 hdif = 2.00e-07 
+rsh = 7.83 rd = 0 rs = 0 
+rsc = 1.5 rdc = 1.5 
// *
// * threshold voltage parameters
// *
+vth0 = -0.402+dvth_p18_rf wvth0 = 1.2675420e-08 pvth0 = -1.2500000e-15+dpvth0_p18_rf 
+k1 = 0.5872390 lk1 = 3.5532110e-09 k2 = 7.0906860e-03 
+k3 = 2.5999999 dvt0 = 0.7194931 dvt1 = 0.2467441 
+dvt2 = 7.8089680e-02 dvt0w = 0.00 dvt1w = 8.0000000e+05 
+dvt2w = 0.00 nlx = 9.0000000e-08 w0 = 0.00 
+k3b = 2.4862001 ngate = 3.1680000e+20 
// *
// * mobility parameters
// *
+vsat = 1.0000000e+05 ua = 2.8500000e-10 lua = 5.5000000e-18 
+pua = -2.0000000e-24 ub = 1.0000000e-18 uc = -4.7700000e-11 
+wuc = 3.1668000e-17 puc = -2.5000000e-24 rdsw = 4.5500000e+02 
+prwb = -0.4000000 prwg = 0.00 wr = 1.0000000 
+u0 = 8.6610000e-03 lu0 = -2.0000000e-11 wu0 = 1.3815350e-10 
+a0 = 1.0000000 keta = 2.0000000e-02 lketa = -8.5000000e-09 
+pketa = 5.0000000e-16 a1 = 0.00 a2 = 0.9900000 
+ags = 0.2000000 b0 = 6.3000000e-08 b1 = 0.00 
// *
// * subthreshold current parameters
// *
+voff = -9.5000000e-02 lvoff = -1.7000000e-09 wvoff = -1.9999999e-09 
+pvoff = -1.0000000e-16 nfactor = 0.9000000 lnfactor = 1.0000000e-07 
+pnfactor = -5.0000000e-15 cit = 0.00 cdsc = 0.00 
+cdscb = 0.00 cdscd = 0.00 eta0 = 4.0000000e-02 
+etab = -2.5000000e-02 dsub = 0.5600000 
// *
// * rout parameters
// *
+pclm = 0.7000000 pdiblc1 = 0.00 pdiblc2 = 7.0000000e-03 
+pdiblcb = 0.00 drout = 0.5600000 pscbe1 = 4.0000000e+08 
+pscbe2 = 1.0000000e-07 pvag = 0.00 delta = 1.0000000e-02 
+alpha0 = 7.0000000e-08 alpha1 = 7.0491700 beta0 = 22.8424000 
+lbeta0 = -7.5000000e-08 
// *
// * temperature effects parameters
// *
+kt1 = -0.2577007 kt2 = -3.0979900e-02 lkt2 = -3.0000000e-09 
+pkt2 = -6.5331750e-16 at = 1.0000000e+04 pat = -1.0000000e-09 
+ute = -1.2703574 ua1 = 5.3866300e-10 wua1 = 1.1000000e-16 
+pua1 = -2.3700001e-24 ub1 = -2.0709999e-18 uc1 = 2.0609721e-11 
+kt1l = -8.0000000e-09 prt = 90.0000000 
// *
// * capacitance parameters
// *
+cj = 0 mj = 0.415 pb = 0.817 
+cjsw = 0 mjsw = 0.489 pbsw = 1 
+cjswg = 0 mjswg = 0.489 pbswg = 1 
+tpb = 0.00153 tpbsw = 0.00117 tpbswg = 0.00117 
+tcj = 0.000876 tcjsw = 0.000745 tcjswg = 0.000745 
+js = 1.66e-07 jsw = 1.2e-13 n = 1.0384 
+xti = 4.5 nqsmod = 0 elm = 5 
+cgdo = cgdo_p18 cgso = cgso_p18 tlevc = 1 
+capmod = 3 xpart = 1 cf = 0.00 
+acde = 0.8505076 moin = 14.95341 noff = 1.431824 
+dlc = -1.5e-09 
+noimod  = 1 flkmod = 1 af = 1.15 kf = 3e-23 
} 
// * junction diode model
model pdio18_rf diode
+is = 1.66e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15 
+n = 1.0135 ns = 1.0135 ik = 4.03e+05 ikp = 2.43e-03 
+bv = 11.0 ibv = 277.78 
+trs = 1.78e-03 eg = 1.16 tnom = 25.0 
+xti = 3.0
+rs = 8.77e-09 
+cjo = 0.00107+dcj_p18_rf 
+cjsw = 5.07e-10+dcjsw_p18_rf
+mj = 0.415 vj = 0.817 mjsw = 0.489 
+vjsw = 1 cta = 0.000876 ctp = 0.000745 
+pta = 0.00153 ptp = 0.00117 tlev = 1 
+tlevc = 1 fc = 0
ends p18_ckt_rf
//*************************
//* 3.3V RF NMOS Subcircuit
//*************************
//* 1=drain, 2=gate, 3=source, 4=bulk
//* lr=gate length, wr=finger width, nf=finger number
subckt n33_ckt_rf (1 2 3 4) 
//* scalable unit parameter
//* euqivalent circuit saclable parameter
parameters lr=0.35u wr=10u nf=2
+rdc_n33_rf      = max(50/(pow(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.7)),1e-3)
+rsc_n33_rf      = max(50/(pow(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.7)),1e-3)
+cgdo_n33_rf     = max((0+dcgdo_n33_rf),0)
+cgso_n33_rf     = max((0+dcgso_n33_rf),0)
//*****************************************
lgate       (2 20)  inductor   l=1p
rgate       (20 21) resistor   r=max((2182.1*lr*1e6+631.05)*pow(nf,(-0.2332*lr*1e6-0.8064))*pow((wr*1e6),((0.028*lr*1e6-0.003)*nf-0.385*lr*1e6-0.7245)),1e-3)
cgd_ext     (20 11) capacitor  c=max((((0.0583*lr*1e6+0.3367)*wr*1e6+(0.2972-0.0222*lr*1e6))*nf+0.4)*1e-15,1e-18)
cgs_ext     (20 31) capacitor  c=max((((2.4814*lr*1e6-0.1584)*log(wr*1e6)+(0.9772*lr*1e6+0.7258))*nf+(3.0576*lr*1e6+1.948))*1e-15,1e-18)
cds_ext     (15 31) capacitor  c=max((3.4-1.8*lr*1e6)*exp((0.047-0.038*lr*1e6)*nf*wr*1e6)*1e-15,1e-18)
rds         (11 15) resistor   r=1m
ldrain      (1 11)  inductor   l=1p
lsource     (3 31)  inductor   l=1p
//*****************************************
djdb (12 11) ndio33_rf area=(nf/2*wr*1e6*(0.8-2*0.07))*1e-12 pj=(1+4.0222e-6*wr*1e6+0.1771/(wr*1e6))*nf*wr
djsb (32 31) ndio33_rf area=(wr*1e6*(0.8-0.07)*2+(nf/2-1)*wr*1e6*(0.8-2*0.07))*1e-12 pj=(1+4.0222e-6*wr*1e6+0.1771/(wr*1e6))*nf*wr
//*****************************************
rsub1      (41  4)  resistor   r=150
rsub2      (41  12) resistor   r=500
rsub3      (41  32) resistor   r=500
//* --------- ideal mos transistor ----------------------
main (11 21 31 41) n33_rf l=lr w=wr m=nf ad = 0 as = 0 pd = 0 ps = 0
// * mos model
model n33_rf bsim3v3 {
1: type=n
// *
// * general parameters
// *
+lmin = 3.3e-7 lmax = 5.2e-7 wmin = 4.8e-7 
+wmax = 1.002e-5 tnom = 25.0 version = 3.2 
+tox = 6.65e-09+dtox_n33_rf toxm = 6.65e-09 xj = 1.6000000e-07 
+nch = 4.3441000e+17 lln = 1.0625758 lwn = 1.0101005 
+wln = 0.9810000 wwn = 0.9060000 lint = 6.3891300e-08 
+ll = -2.3305548e-15 lw = -2.4634918e-15 lwl = 2.6243002e-24 
+wint = 3.5850000e-08 wl = -1.8902563e-15 ww = -1.3000000e-14 
+wwl = -1.3027796e-20 mobmod = 1 binunit = 2 
+xl = 1e-8+dxl_n33_rf xw = 0.00+dxw_n33_rf dwg = -3.9100000e-09 
+dwb = 3.2000000e-09 
// * diode parameters
+dskip = no ldif = 6.50e-08 hdif = 2.05e-07 
+rsh = 7.08 rd = 0 rs = 0 
+rsc = rsc_n33_rf rdc = rdc_n33_rf 
// *
// * threshold voltage parameters
// *
+vth0 = 0.695+dvth_n33_rf lvth0 = 4.0100000e-10 wvth0 = 1.0200000e-08 
+pvth0 = 8.0000000e-16+dpvth0_n33_rf k1 = 0.8451000 lk1 = 5.8182560e-10 
+wk1 = -6.2456240e-09 pk1 = 1.9938927e-15 k2 = 4.4575000e-02 
+k3 = -3.8500000 dvt0 = 9.4991400 ldvt0 = 8.0839730e-09 
+dvt1 = 0.6300000 ldvt1 = 5.5000000e-08 dvt2 = -0.1450000 
+dvt0w = 0.00 dvt1w = 0.1057000 dvt2w = 0.00 
+nlx = 2.0274594e-07 lnlx = -2.8608589e-14 w0 = 0.00 
+k3b = 0.5669292 ngate = 2.6812141e+21 
// *
// * mobility parameters
// *
+vsat = 8.5000000e+04 lvsat = -1.7300000e-03 pvsat = 1.2000000e-10 
+ua = -8.6001130e-10 ub = 2.3000001e-18 uc = 1.3100000e-10 
+puc = 5.0000000e-25 rdsw = 2.4208382e+02 prwb = -8.5000000e-02 
+prwg = 3.8000000e-02 wr = 1.0000000 u0 = 3.5000000e-02 
+lu0 = 5.0000000e-10 a0 = 1.0200000 la0 = -1.2000000e-07 
+keta = 0.00 lketa = -1.4000000e-08 wketa = -1.9999999e-09 
+pketa = 1.0000000e-15 a1 = 0.00 a2 = 0.9900000 
+ags = 0.1700000 b0 = 1.0000000e-08 b1 = 0.00 
// *
// * subthreshold current parameters
// *
+voff = -0.1200000 nfactor = 1.1000000 lnfactor = 4.0000000e-08 
+pnfactor = -1.4000000e-14 cit = 1.0000000e-04 cdsc = 5.0000000e-04 
+cdscb = 0.00 cdscd = 0.00 eta0 = 4.0000000e-02 
+peta0 = 3.0000001e-16 etab = -0.1000000 dsub = 0.6000000 
// *
// * rout parameters
// *
+pclm = 0.8000000 lpclm = 5.0000000e-08 ppclm = 8.0000000e-15 
+pdiblc1 = 9.0000000e-02 pdiblc2 = 1.6000000e-03 ppdiblc2 = -7.0000000e-17 
+pdiblcb = 0.00 drout = 0.5987002 pscbe1 = 3.4000000e+08 
+lpscbe1 = 13.0000000 pscbe2 = 3.8000000e-06 pvag = 0.00 
+delta = 1.0000000e-02 alpha0 = -4.4760000e-08 alpha1 = 0.8998877 
+beta0 = 18.8771250 lbeta0 = -5.7118000e-07 
// *
// * temperature effects parameters
// *
+kt1 = -0.3250000 pkt1 = -2.3708420e-15 kt2 = -3.6844640e-02 
+at = 2.2000000e+04 ute = -1.4100000 ua1 = 2.0599999e-09 
+wua1 = -1.2600000e-16 pua1 = -1.0000000e-24 ub1 = -2.5000000e-18 
+wub1 = 1.1000000e-25 uc1 = -1.1000000e-10 luc1 = 1.6999999e-17 
+kt1l = -5.0000000e-09 prt = 40.0000000 
// *
// *
// * capacitance parameters
// *
+cj = 0 mj = 0.321 pb = 0.708 
+cjsw = 0 mjsw = 0.447 pbsw = 1 
+cjswg = 0 mjswg = 0.447 pbswg = 1 
+tpb = 0.00166 tpbsw = 0.00162 tpbswg = 0.00162 
+tcj = 0.000897 tcjsw = 0.000695 tcjswg = 0.000695 
+js = 3.65e-07 jsw = 3.0e-13 n = 1.04 
+xti = 3.9 nqsmod = 0 elm = 5 
+cgdo = cgdo_n33_rf cgso = cgso_n33_rf tlevc = 1 
+capmod = 3 xpart = 1 cf = 0.00 
+acde = 0.45 moin = 24 noff = 2.3177 
+dlc = 6.50e-08 
+noimod  = 1 flkmod = 1 af = 1 kf = 3e-23 
}
// * junction diode model
model ndio33_rf diode
+is = 3.65e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15 
+n = 1.0203 ns = 1.0203 rs = 8.84e-09 ik = 1.33e+05 ikp = 3.64e-04 
+bv = 11.0 ibv = 277.78 
+trs = 1.07e-03 eg = 1.16 tnom = 25.0 
+xti = 3.0 cjo = 0.000845+dcj_n33_rf mj = 0.321 
+vj = 0.708 cjsw = 3.41e-10+dcjsw_n33_rf mjsw = 0.447 
+vjsw = 1 cta = 0.000897 ctp = 0.000695 
+pta = 0.00166 ptp = 0.00162 tlev = 1 
+tlevc = 1 fc = 0 
ends n33_ckt_rf
//***************************
//* 3.3V RF DNWMOS Subcircuit
//***************************
//* 1=drain, 2=gate, 3=source, 4=bulk, 5=DNW
//* lr=gate length, wr=finger width, nf=finger number, laddr=DNW diode add length, waddr=DNW diode add width
subckt dnw33_ckt_rf (1 2 3 4 5) 
//* scalable unit parameter
//* euqivalent circuit saclable parameter
parameters lr=0.35u wr=10u nf=2 laddr=10u waddr=10u
+rdc_n33_rf      = max(50/(pow(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.7)),1e-3)
+rsc_n33_rf      = max(50/(pow(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.7)),1e-3)
+cgdo_n33_rf     = max((0+dcgdo_n33_rf),0)
+cgso_n33_rf     = max((0+dcgso_n33_rf),0)
//*****************************************
lgate       (2 20)  inductor   l=1p
rgate       (20 21) resistor   r=max((2182.1*lr*1e6+631.05)*pow(nf,(-0.2332*lr*1e6-0.8064))*pow((wr*1e6),((0.028*lr*1e6-0.003)*nf-0.385*lr*1e6-0.7245)),1e-3)
cgd_ext     (20 11) capacitor  c=max((((0.0583*lr*1e6+0.3367)*wr*1e6+(0.2972-0.0222*lr*1e6))*nf+0.4)*1e-15,1e-18)
cgs_ext     (20 31) capacitor  c=max((((2.4814*lr*1e6-0.1584)*log(wr*1e6)+(0.9772*lr*1e6+0.7258))*nf+(3.0576*lr*1e6+1.948))*1e-15,1e-18)
cds_ext     (15 31) capacitor  c=max((3.4-1.8*lr*1e6)*exp((0.047-0.038*lr*1e6)*nf*wr*1e6)*1e-15,1e-18)
rds         (11 15) resistor   r=1m
ldrain      (1 11)  inductor   l=1p
lsource     (3 31)  inductor   l=1p
//*****************************************
djdb (12 11) ndio33_rf area=(nf/2*wr*1e6*(0.8-2*0.07))*1e-12 pj=(1+4.0222e-6*wr*1e6+0.1771/(wr*1e6))*nf*wr
djsb (32 31) ndio33_rf area=(wr*1e6*(0.8-0.07)*2+(nf/2-1)*wr*1e6*(0.8-2*0.07))*1e-12 pj=(1+4.0222e-6*wr*1e6+0.1771/(wr*1e6))*nf*wr
djdnw (4 5) diobpw_rf area=(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+2*laddr)*(wr+2*waddr) pj=2*(2*0.8*1e-6+lr*nf+0.8*1e-6*(nf-1)+wr+2*(laddr+waddr))
//*****************************************
rsub1      (41  4)  resistor   r=150
rsub2      (41  12) resistor   r=500
rsub3      (41  32) resistor   r=500
//* --------- ideal mos transistor ----------------------
main (11 21 31 41) dnw33_rf l=lr w=wr m=nf ad = 0 as = 0 pd = 0 ps = 0
// * mos model
model dnw33_rf bsim3v3 {
1: type=n
// *
// * general parameters
// *
+lmin = 3.3e-7 lmax = 5.2e-7 wmin = 4.8e-7 
+wmax = 1.002e-5 tnom = 25.0 version = 3.2 
+tox = 6.65e-09+dtox_n33_rf toxm = 6.65e-09 xj = 1.6000000e-07 
+nch = 4.3441000e+17 lln = 1.0625758 lwn = 1.0101005 
+wln = 0.9810000 wwn = 0.9060000 lint = 6.3891300e-08 
+ll = -2.3305548e-15 lw = -2.4634918e-15 lwl = 2.6243002e-24 
+wint = 3.5850000e-08 wl = -1.8902563e-15 ww = -1.3000000e-14 
+wwl = -1.3027796e-20 mobmod = 1 binunit = 2 
+xl = 1e-8+dxl_n33_rf xw = 0.00+dxw_n33_rf dwg = -3.9100000e-09 
+dwb = 3.2000000e-09 
// * diode parameters
+dskip = no ldif = 6.50e-08 hdif = 2.05e-07 
+rsh = 7.08 rd = 0 rs = 0 
+rsc = rsc_n33_rf rdc = rdc_n33_rf 
// *
// * threshold voltage parameters
// *
+vth0 = 0.695+dvth_n33_rf lvth0 = 4.0100000e-10 wvth0 = 1.0200000e-08 
+pvth0 = 8.0000000e-16+dpvth0_n33_rf k1 = 0.8451000 lk1 = 5.8182560e-10 
+wk1 = -6.2456240e-09 pk1 = 1.9938927e-15 k2 = 4.4575000e-02 
+k3 = -3.8500000 dvt0 = 9.4991400 ldvt0 = 8.0839730e-09 
+dvt1 = 0.6300000 ldvt1 = 5.5000000e-08 dvt2 = -0.1450000 
+dvt0w = 0.00 dvt1w = 0.1057000 dvt2w = 0.00 
+nlx = 2.0274594e-07 lnlx = -2.8608589e-14 w0 = 0.00 
+k3b = 0.5669292 ngate = 2.6812141e+21 
// *
// * mobility parameters
// *
+vsat = 8.5000000e+04 lvsat = -1.7300000e-03 pvsat = 1.2000000e-10 
+ua = -8.6001130e-10 ub = 2.3000001e-18 uc = 1.3100000e-10 
+puc = 5.0000000e-25 rdsw = 2.4208382e+02 prwb = -8.5000000e-02 
+prwg = 3.8000000e-02 wr = 1.0000000 u0 = 3.5000000e-02 
+lu0 = 5.0000000e-10 a0 = 1.0200000 la0 = -1.2000000e-07 
+keta = 0.00 lketa = -1.4000000e-08 wketa = -1.9999999e-09 
+pketa = 1.0000000e-15 a1 = 0.00 a2 = 0.9900000 
+ags = 0.1700000 b0 = 1.0000000e-08 b1 = 0.00 
// *
// * subthreshold current parameters
// *
+voff = -0.1200000 nfactor = 1.1000000 lnfactor = 4.0000000e-08 
+pnfactor = -1.4000000e-14 cit = 1.0000000e-04 cdsc = 5.0000000e-04 
+cdscb = 0.00 cdscd = 0.00 eta0 = 4.0000000e-02 
+peta0 = 3.0000001e-16 etab = -0.1000000 dsub = 0.6000000 
// *
// * rout parameters
// *
+pclm = 0.8000000 lpclm = 5.0000000e-08 ppclm = 8.0000000e-15 
+pdiblc1 = 9.0000000e-02 pdiblc2 = 1.6000000e-03 ppdiblc2 = -7.0000000e-17 
+pdiblcb = 0.00 drout = 0.5987002 pscbe1 = 3.4000000e+08 
+lpscbe1 = 13.0000000 pscbe2 = 3.8000000e-06 pvag = 0.00 
+delta = 1.0000000e-02 alpha0 = -4.4760000e-08 alpha1 = 0.8998877 
+beta0 = 18.8771250 lbeta0 = -5.7118000e-07 
// *
// * temperature effects parameters
// *
+kt1 = -0.3250000 pkt1 = -2.3708420e-15 kt2 = -3.6844640e-02 
+at = 2.2000000e+04 ute = -1.4100000 ua1 = 2.0599999e-09 
+wua1 = -1.2600000e-16 pua1 = -1.0000000e-24 ub1 = -2.5000000e-18 
+wub1 = 1.1000000e-25 uc1 = -1.1000000e-10 luc1 = 1.6999999e-17 
+kt1l = -5.0000000e-09 prt = 40.0000000 
// *
// *
// * capacitance parameters
// *
+cj = 0 mj = 0.321 pb = 0.708 
+cjsw = 0 mjsw = 0.447 pbsw = 1 
+cjswg = 0 mjswg = 0.447 pbswg = 1 
+tpb = 0.00166 tpbsw = 0.00162 tpbswg = 0.00162 
+tcj = 0.000897 tcjsw = 0.000695 tcjswg = 0.000695 
+js = 3.65e-07 jsw = 3.0e-13 n = 1.04 
+xti = 3.9 nqsmod = 0 elm = 5 
+cgdo = cgdo_n33_rf cgso = cgso_n33_rf tlevc = 1 
+capmod = 3 xpart = 1 cf = 0.00 
+acde = 0.45 moin = 24 noff = 2.3177 
+dlc = 6.50e-08 
+noimod  = 1 flkmod = 1 af = 1 kf = 3e-23 
}
// * junction diode model
model ndio33_rf diode
+is = 3.65e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15 
+n = 1.0203 ns = 1.0203 rs = 8.84e-09 ik = 1.33e+05 ikp = 3.64e-04 
+bv = 11.0 ibv = 277.78 
+trs = 1.07e-03 eg = 1.16 tnom = 25.0 
+xti = 3.0 cjo = 0.000845+dcj_n33_rf mj = 0.321 
+vj = 0.708 cjsw = 3.41e-10+dcjsw_n33_rf mjsw = 0.447 
+vjsw = 1 cta = 0.000897 ctp = 0.000695 
+pta = 0.00166 ptp = 0.00162 tlev = 1 
+tlevc = 1 fc = 0 
// * DNW junction diode model
model diobpw_rf diode
+level = 1 is = 1.50e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1.00e-15 
+n = 1.0213 ns = 1.0213 rs = 2.51e-08 ik = 2.40e+05 ikp = 1.60E-03 
+bv = 15.0 ibv = 1.04e+02 
+trs = 1.77e-03 cta = 0.0012 ctp = 0.00107 
+eg = 1.16 tnom = 25.0 pta = 0.0019 
+ptp = 0.00193 xti = 3.0 cjo = 0.000536 
+mj = 0.343 vj = 0.693 cjsw = 3.22e-10 
+mjsw = 0.361 vjsw = 0.715 tlev = 1 
+tlevc = 1 area = 9.6e-9 perim = 4e-4 
+fc = 0 
ends dnw33_ckt_rf
//*************************
//* 3.3V RF PMOS Subcircuit
//*************************
//* 1=drain, 2=gate, 3=source, 4=bulk
//* lr=gate length, wr=finger width, nf=finger number
subckt p33_ckt_rf (1 2 3 4) 
//* scalable unit parameter
//* euqivalent circuit saclable parameter
parameters lr=0.3u wr=10u nf=2
+rdc_p33_rf      = max(81.5/(pow(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.95)),1e-3)
+rsc_p33_rf      = max(81.5/(pow(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.95)),1e-3)
+cgdo_p33_rf     = max((0+dcgdo_p33_rf),0)
+cgso_p33_rf     = max((0+dcgso_p33_rf),0)
//*****************************************
lgate       (2 20)  inductor   l=1p
rgate       (20 21) resistor   r=max((6345.5*lr*1e6+389.25)*pow(nf,(0.303*lr*1e6-1.1215))*pow((wr*1e6),(-0.6785*lr*1e6-0.4944)),1e-3)
cgd_ext     (20 11) capacitor  c=max(((0.1595*lr*1e6+0.2682)*wr*1e6*nf+(0.255+0.058*lr*1e6)*nf+0.8393-1.1375*lr*1e6)*1e-15,1e-18)
cgs_ext     (20 31) capacitor  c=max((((0.3785-0.0165*lr*1e6)*wr*1e6+(0.9772*lr*1e6+0.1732))*nf+4)*1e-15,1e-18)
cds_ext     (15 31) capacitor  c=max(((0.8638-0.8045*lr*1e6)*wr*1e6+(1.9425*lr*1e6-0.7838))*nf*1e-15,1e-18)
rds         (11 15) resistor   r=80.2
ldrain      (1 11)  inductor   l=1p
lsource     (3 31)  inductor   l=1p
//*****************************************
djdb (11 12) pdio33_rf area=(nf/2*wr*1e6*(0.8-2*0.07))*1e-12 pj=(1-6.0826e-6*wr*1e6+0.1854/wr*1e6)*nf*wr
djsb (31 32) pdio33_rf area=(wr*1e6*(0.8-0.07)*2+(nf/2-1)*wr*1e6*(0.8-2*0.07))*1e-12 pj=(1-6.0826e-6*wr*1e6+0.1854/wr*1e6)*nf*wr
//*****************************************
rsub1      (41  4)  resistor   r=10
rsub2      (41  12) resistor   r=50000
rsub3      (41  32) resistor   r=50000
//* --------- ideal mos transistor ----------------------
main (11 21 31 41) p33_rf l=lr w=wr m=nf ad = 0 as = 0 pd = 0 ps = 0
// * mos model
model p33_rf bsim3v3 {
1: type=p
// *
// * general parameters
// *
+lmin = 2.8e-7 lmax = 5.2e-7 wmin = 4.8e-7 
+wmax = 1.002e-5 tnom = 25.0 version = 3.2 
+tox = 6.62e-09+dtox_p33_rf toxm = 6.62e-09 xj = 1.7000001e-07 
+nch = 5.4852000e+17 lln = 1.0471729 lwn = 0.9530895 
+wln = 1.0257638 wwn = 0.9617700 lint = 3.5000000e-08 
+ll = 5.5000000e-15 lw = -4.7160380e-14 lwl = 7.0054450e-22 
+wint = 1.3000000e-08 wl = -3.1491245e-14 ww = 2.3000000e-15 
+wwl = -2.4167156e-22 mobmod = 1 binunit = 2 
+xl = -1.70e-08+dxl_p33_rf xw = 0.00+dxw_p33_rf dwg = 0.00 
+dwb = 8.6000000e-09 
// * diode parameters
+dskip = no ldif = 6.50e-08 hdif = 2.05e-07 
+rsh = 9.8 rd = 0 rs = 0 
+rsc = rsc_p33_rf rdc = rdc_p33_rf 
// *
// * threshold voltage parameters
// *
+vth0 = -0.672+dvth_p33_rf wvth0 = 4.0000000e-09 pvth0 = 6.0000000e-15+dpvth0_p33_rf 
+k1 = 0.9145741 pk1 = -1.7000000e-14 k2 = 4.1276220e-02 
+k3 = 0.1293833 dvt0 = 1.8000000 dvt1 = 0.7100000 
+dvt2 = -7.0000000e-02 dvt0w = 0.00 dvt1w = 0.00 
+dvt2w = 0.00 nlx = 1.2000000e-08 w0 = 1.0021131e-09 
+k3b = 0.4000000 ngate = 1.1600000e+20 
// *
// * mobility parameters
// *
+vsat = 8.5500000e+04 pvsat = -5.8000000e-09 ua = 3.1500000e-10 
+lua = 1.5000001e-17 wua = -1.6763224e-16 pua = -1.1000000e-23 
+ub = 1.0444180e-18 lub = -7.0000000e-27 uc = -3.5000000e-11 
+luc = 4.0000000e-18 puc = 5.0000000e-24 rdsw = 9.5000000e+02 
+prwb = 0.00 prwg = 6.3755660e-03 wr = 1.0000000 
+u0 = 9.2500000e-03 lu0 = -4.1500680e-10 wu0 = -1.7001526e-12 
+pu0 = -3.7999640e-16 a0 = 0.8500000 keta = 1.5000000e-02 
+lketa = -1.0000000e-08 wketa = 1.0000000e-09 pketa = -6.0000000e-15 
+a1 = 0.00 a2 = 0.9900000 ags = 4.0000000e-02 
+b0 = 4.6000000e-08 b1 = 0.00 
// *
// * subthreshold current parameters
// *
+voff = -0.1000000 lvoff = 1.8000000e-09 pvoff = -2.9999999e-15 
+nfactor = 1.1000000 pnfactor = -4.0000000e-14 cit = 1.9999999e-04 
+cdsc = 4.5263850e-05 cdscb = 0.00 cdscd = 0.00 
+eta0 = 5.0000000e-03 peta0 = 7.0000000e-15 etab = -1.5000000e-02 
+petab = -2.0000000e-15 dsub = 0.5800000 
// *
// * rout parameters
// *
+pclm = 0.6000000 ppclm = 1.3000000e-13 pdiblc1 = 6.0000000e-03 
+pdiblc2 = 2.5000001e-04 wpdiblc2 = 8.0000000e-11 pdiblcb = 0.00 
+drout = 0.5600000 pscbe1 = 3.3000000e+08 ppscbe1 = -7.0000000e-06 
+pscbe2 = 2.0000000e-07 pvag = 0.00 delta = 8.0000000e-03 
+pdelta = 4.0000000e-16 alpha0 = 1.3410400e-06 alpha1 = 5.6136910e-02 
+beta0 = 27.5998000 
// *
// * temperature effects parameters
// *
+kt1 = -0.3840900 wkt1 = -9.4333370e-10 pkt1 = 4.9999980e-15 
+kt2 = -4.1563480e-02 at = -2.0000000e+03 pat = -7.5000000e-09 
+ute = -1.3236057 ua1 = 3.0000002e-10 wua1 = 8.0000000e-18 
+pua1 = 1.0000000e-23 ub1 = -2.0704662e-18 wub1 = 1.4000000e-25 
+uc1 = -5.0000000e-11 kt1l = -6.0000000e-09 prt = 1.3000000e+02 
// *
// * capacitance parameters
// *
+cj = 0 mj = 0.401 pb = 0.807 
+cjsw = 0 mjsw = 0.45 pbsw = 1 
+cjswg = 0 mjswg = 0.45 pbswg = 1 
+tpb = 0.00157 tpbsw = 0.00137 tpbswg = 0.00137 
+tcj = 0.000883 tcjsw = 0.000709 tcjswg = 0.000709 
+js = 1.68e-07 jsw = 4.0e-13 n = 1.07 
+xti = 3.0 nqsmod = 0 elm = 5 
+cgdo = cgdo_p33_rf cgso = cgdo_p33_rf tlevc = 1 
+capmod = 3 xpart = 1 cf = 0.00 
+acde = 0.55 moin = 15 noff = 0.565 
+dlc = 7.0e-09 dwc = 6.0e-8 
+noimod  = 1 flkmod = 1 af = 1.02 kf = 3e-23
} 
// * junction diode model
model pdio33_rf diode
+is = 1.68e-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15 
+n = 1.0143 ns = 1.0143 rs = 9.23e-09 ik = 4.07e+05 ikp = 2.42e-03 
+bv = 11.0 ibv = 277.78 
+trs = 1.24e-03 eg = 1.16 tnom = 25.0 
+xti = 3.0 cjo = 0.00101+dcj_p33_rf mj = 0.401 
+vj = 0.807 cjsw = 3.19e-10+dcjsw_p33_rf mjsw = 0.45 
+vjsw = 1 cta = 0.000883 ctp = 0.000709 
+pta = 0.00157 ptp = 0.00137 tlev = 1 
+tlevc = 1 fc = 0 
ends p33_ckt_rf
//*
