* SPICE NETLIST
***************************************

.SUBCKT And_Gate VIN_B VIN_A VDD GND VOUT
** N=7 EP=5 IP=0 FDC=6
M0 6 VIN_A 7 GND NM L=1.8e-07 W=2.2e-07 $X=1890 $Y=-4485 $D=0
M1 GND VIN_B 6 GND NM L=1.8e-07 W=2.2e-07 $X=2690 $Y=-4485 $D=0
M2 VOUT 7 GND GND NM L=1.8e-07 W=2.2e-07 $X=3490 $Y=-4485 $D=0
M3 7 VIN_A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1890 $Y=-2095 $D=4
M4 VDD VIN_B 7 VDD PM L=1.8e-07 W=4.4e-07 $X=2610 $Y=-2095 $D=4
M5 VOUT 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3330 $Y=-2095 $D=4
.ENDS
***************************************
.SUBCKT AND_5 A B C VDD GND E D OUT
** N=13 EP=8 IP=10 FDC=20
M0 5 A 9 GND NM L=1.8e-07 W=2.2e-07 $X=2675 $Y=-19050 $D=0
M1 6 B 5 GND NM L=1.8e-07 W=2.2e-07 $X=3475 $Y=-19050 $D=0
M2 GND C 6 GND NM L=1.8e-07 W=2.2e-07 $X=4275 $Y=-19050 $D=0
M3 4 9 GND GND NM L=1.8e-07 W=2.2e-07 $X=5075 $Y=-19050 $D=0
M4 VDD A 9 VDD PM L=1.8e-07 W=4.4e-07 $X=2755 $Y=-16660 $D=4
M5 9 B VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3475 $Y=-16660 $D=4
M6 VDD C 9 VDD PM L=1.8e-07 W=4.4e-07 $X=4195 $Y=-16660 $D=4
M7 4 9 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=4915 $Y=-16660 $D=4
X8 E D VDD GND 10 And_Gate $T=4715 -14565 0 0 $X=5695 $Y=-20190
X9 10 4 VDD GND OUT And_Gate $T=7865 -14565 0 0 $X=8845 $Y=-20190
.ENDS
***************************************
