* SPICE NETLIST
***************************************

.SUBCKT n18_2 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT RAM_v1 WL Q BL GND VDD
** N=7 EP=5 IP=20 FDC=8
X0 GND 7 6 WL n18_2 $T=2520 -3795 0 0 $X=1820 $Y=-4935
X1 GND Q BL WL n18_2 $T=7180 -3795 0 0 $X=6480 $Y=-4935
X2 6 GND VDD Q inv $T=7305 -8020 0 0 $X=3190 $Y=-4935
X3 Q GND VDD 6 inv $T=8805 -8020 0 0 $X=4690 $Y=-4935
X4 BL GND VDD 7 inv $T=11965 -8020 0 0 $X=7850 $Y=-4935
.ENDS
***************************************
.SUBCKT 12_RAM_v1 WL Q<11> B<11> Q<10> B<10> Q<9> B<9> Q<8> B<8> Q<7> B<7> Q<6> B<6> Q<5> B<5> Q<4> B<4> Q<3> B<3> Q<2>
+ B<2> Q<1> B<1> Q<0> B<0> GND VDD
** N=27 EP=27 IP=60 FDC=96
X0 WL Q<11> B<11> GND VDD RAM_v1 $T=1705 -46690 0 0 $X=3525 $Y=-51665
X1 WL Q<10> B<10> GND VDD RAM_v1 $T=1705 -42535 0 0 $X=3525 $Y=-47510
X2 WL Q<9> B<9> GND VDD RAM_v1 $T=1705 -38385 0 0 $X=3525 $Y=-43360
X3 WL Q<8> B<8> GND VDD RAM_v1 $T=1705 -34220 0 0 $X=3525 $Y=-39195
X4 WL Q<7> B<7> GND VDD RAM_v1 $T=1705 -30055 0 0 $X=3525 $Y=-35030
X5 WL Q<6> B<6> GND VDD RAM_v1 $T=1705 -25900 0 0 $X=3525 $Y=-30875
X6 WL Q<5> B<5> GND VDD RAM_v1 $T=1705 -21750 0 0 $X=3525 $Y=-26725
X7 WL Q<4> B<4> GND VDD RAM_v1 $T=1705 -17585 0 0 $X=3525 $Y=-22560
X8 WL Q<3> B<3> GND VDD RAM_v1 $T=1705 -13430 0 0 $X=3525 $Y=-18405
X9 WL Q<2> B<2> GND VDD RAM_v1 $T=1705 -9280 0 0 $X=3525 $Y=-14255
X10 WL Q<1> B<1> GND VDD RAM_v1 $T=1705 -5125 0 0 $X=3525 $Y=-10100
X11 WL Q<0> B<0> GND VDD RAM_v1 $T=1705 -975 0 0 $X=3525 $Y=-5950
.ENDS
***************************************
