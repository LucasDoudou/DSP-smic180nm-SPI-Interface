//* 
//* No part of this file can be released without the consent of SMIC.
//*
//******************************************************************************************
//* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.6
//*
//* Release date       : 07/02/2007
//*
//* Simulation tool    : Cadence spectre V6.0
//*
//*
//*  MIM Capacitor   :
//*
//*        *--------------------------------* 
//*        |  1fF/um^2 subckt  |  mim1__rf  |
//*        *--------------------------------*
simulator lang=spectre  insensitive=yes
//*******************************
//* 0.18um 1fF/um^2 MIM Capacitor
//*******************************
//* 1=port1, 2=port2
subckt mim1_rf (1 2)
//* mim capacitor scalable model parameters
parameters lr=10 wr=10
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1465+6.59474/(lr*wr*1E12)+215.51267/((lr*wr*1E12)*(lr*wr*1E12)))*1E-9, 1E-13)
cf    (22 2)  mim1       l=lr w=wr
rs    (11 22) resistor   r=max(0.24417+185.93086/(lr*wr*1E12), 1E-6)
rsub1 (10 0)  resistor   r=max(3.0E+04-2.0*lr*wr*1E12, 1E-3)
csub1 (10 0)  capacitor  c=max((0.08*lr*1E6)*1E-15, 1E-18)
cox1  (1 10)  capacitor  c=max((2.5E-03*lr*wr*1E12)*1E-15, 1E-18)
rsub2 (20 0)  resistor   r=max(4.88E+03-0.6495*lr*wr*1E12, 1E-3)
csub2 (20 0)  capacitor  c=max((0.1*lr*1E6)*1E-15, 1E-18)
cox2  (2 20)  capacitor  c=max((6.38E-03*lr*wr*1E12)*1E-15, 1E-18)
ends mim1_rf
//*********************
model mim1 capacitor
+coeffs = [-3.411E-5 -1.489E-5]
+tc1 = -3.482E-05  tnom = 25
+cj = 1E-03+dmim1_rf
