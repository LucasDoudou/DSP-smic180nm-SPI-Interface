* SPICE NETLIST
***************************************

.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Cobar CI B A GND VDD CO_
** N=10 EP=6 IP=24 FDC=10
M0 7 CI CO_ GND NM L=1.8e-07 W=4.4e-07 $X=8000 $Y=-13525 $D=0
M1 6 CI CO_ VDD PM L=1.8e-07 W=8.8e-07 $X=8000 $Y=-9500 $D=4
X2 VDD 6 VDD 6 B A p18_0 $T=9495 -9500 0 0 $X=8585 $Y=-9930
X3 VDD CO_ 10 VDD B A p18_0 $T=11715 -9500 0 0 $X=10805 $Y=-9930
X4 GND GND 7 B A n18_2 $T=9495 -13525 0 0 $X=8835 $Y=-14655
X5 GND CO_ 9 B A n18_2 $T=11715 -13525 0 0 $X=11055 $Y=-14655
.ENDS
***************************************
