* SPICE NETLIST
***************************************

.SUBCKT And_Gate VIN_B VIN_A VDD GND VOUT
** N=7 EP=5 IP=0 FDC=6
M0 6 VIN_A 7 GND NM L=1.8e-07 W=2.2e-07 $X=1890 $Y=-4485 $D=0
M1 GND VIN_B 6 GND NM L=1.8e-07 W=2.2e-07 $X=2690 $Y=-4485 $D=0
M2 VOUT 7 GND GND NM L=1.8e-07 W=2.2e-07 $X=3490 $Y=-4485 $D=0
M3 7 VIN_A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1890 $Y=-2095 $D=4
M4 VDD VIN_B 7 VDD PM L=1.8e-07 W=4.4e-07 $X=2610 $Y=-2095 $D=4
M5 VOUT 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3330 $Y=-2095 $D=4
.ENDS
***************************************
.SUBCKT 6_AND_test Y<0> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND Z<0> A<0> A<1> A<2> A<3> A<4>
** N=15 EP=15 IP=30 FDC=36
X0 X<0> Y<0> VDD GND Z<0> And_Gate $T=2375 -2105 0 0 $X=3355 $Y=-7730
X1 X<1> Y<0> VDD GND A<0> And_Gate $T=5555 -2105 0 0 $X=6535 $Y=-7730
X2 X<2> Y<0> VDD GND A<1> And_Gate $T=8735 -2105 0 0 $X=9715 $Y=-7730
X3 X<3> Y<0> VDD GND A<2> And_Gate $T=11915 -2105 0 0 $X=12895 $Y=-7730
X4 X<4> Y<0> VDD GND A<3> And_Gate $T=15095 -2105 0 0 $X=16075 $Y=-7730
X5 X<5> Y<0> VDD GND A<4> And_Gate $T=18275 -2105 0 0 $X=19255 $Y=-7730
.ENDS
***************************************
.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT 6_FA_v3 S<0> S<1> S<2> S<3> S<4> S<5> S<6> A<0> B<0> GND A<1> B<1> A<2> B<2> A<3> B<3> A<4> B<4> A<5> B<5>
+ VDD
** N=38 EP=21 IP=78 FDC=168
X0 33 GND VDD S<0> 22 29 ICV_1 $T=11635 -18360 0 0 $X=7520 $Y=-15275
X1 34 GND VDD S<1> 23 30 ICV_1 $T=11635 -10670 0 0 $X=7520 $Y=-7585
X2 35 GND VDD S<2> 24 31 ICV_1 $T=11635 -2795 0 0 $X=7520 $Y=290
X3 36 GND VDD S<3> 25 28 ICV_1 $T=11635 4895 0 0 $X=7520 $Y=7980
X4 37 GND VDD S<4> 26 32 ICV_1 $T=11635 12720 0 0 $X=7520 $Y=15805
X5 38 GND VDD S<5> 27 S<6> ICV_1 $T=11635 20410 0 0 $X=7520 $Y=23495
X6 GND A<0> B<0> 22 GND VDD 33 Full_Adder_Sum $T=-17990 4290 0 0 $X=-7550 $Y=-15275
X7 29 A<1> B<1> 23 GND VDD 34 Full_Adder_Sum $T=-17990 11980 0 0 $X=-7550 $Y=-7585
X8 30 A<2> B<2> 24 GND VDD 35 Full_Adder_Sum $T=-17990 19855 0 0 $X=-7550 $Y=290
X9 31 A<3> B<3> 25 GND VDD 36 Full_Adder_Sum $T=-17990 27545 0 0 $X=-7550 $Y=7980
X10 28 A<4> B<4> 26 GND VDD 37 Full_Adder_Sum $T=-17990 35370 0 0 $X=-7550 $Y=15805
X11 32 A<5> B<5> 27 GND VDD 38 Full_Adder_Sum $T=-17990 43060 0 0 $X=-7550 $Y=23495
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=12
X0 1 3 4 5 6 And_Gate $T=0 0 0 0 $X=980 $Y=-5625
X1 2 3 4 5 7 And_Gate $T=3180 0 0 0 $X=4160 $Y=-5625
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=24
X0 1 2 7 6 5 8 9 ICV_2 $T=0 0 0 0 $X=980 $Y=-5625
X1 3 4 10 6 5 11 12 ICV_2 $T=6360 0 0 0 $X=7340 $Y=-5625
.ENDS
***************************************
.SUBCKT 5_6_Multiplier X<0> X<1> X<2> X<3> X<4> X<5> Y<1> Y<0> Z<0> Z<1> GND Y<3> Y<4> Y<2> Z<5> Z<6> Z<7> Z<8> Z<9> Z<10>
+ VDD Z<2> Z<3> Z<4>
** N=88 EP=24 IP=222 FDC=852
X0 Y<2> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 52 53 54 55 56 57 6_AND_test $T=51110 -22420 0 0 $X=54270 $Y=-30150
X1 Y<3> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 59 60 61 62 63 64 6_AND_test $T=75810 -22420 0 0 $X=78970 $Y=-30150
X2 Y<4> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 66 67 68 69 70 71 6_AND_test $T=100535 -22420 0 0 $X=103695 $Y=-30150
X3 80 GND VDD Z<1> 39 48 ICV_1 $T=48685 -77935 0 0 $X=44570 $Y=-74850
X4 81 GND VDD 15 40 49 ICV_1 $T=48685 -70245 0 0 $X=44570 $Y=-67160
X5 82 GND VDD 16 41 50 ICV_1 $T=48685 -62370 0 0 $X=44570 $Y=-59285
X6 83 GND VDD 18 42 47 ICV_1 $T=48685 -54680 0 0 $X=44570 $Y=-51595
X7 84 GND VDD 14 43 51 ICV_1 $T=48685 -46855 0 0 $X=44570 $Y=-43770
X8 85 GND VDD 17 44 13 ICV_1 $T=48685 -39165 0 0 $X=44570 $Y=-36080
X9 GND 34 7 39 GND VDD 80 Full_Adder_Sum $T=19060 -55285 0 0 $X=29500 $Y=-74850
X10 48 35 8 40 GND VDD 81 Full_Adder_Sum $T=19060 -47595 0 0 $X=29500 $Y=-67160
X11 49 36 9 41 GND VDD 82 Full_Adder_Sum $T=19060 -39720 0 0 $X=29500 $Y=-59285
X12 50 37 10 42 GND VDD 83 Full_Adder_Sum $T=19060 -32030 0 0 $X=29500 $Y=-51595
X13 47 38 11 43 GND VDD 84 Full_Adder_Sum $T=19060 -24205 0 0 $X=29500 $Y=-43770
X14 51 GND 12 44 GND VDD 85 Full_Adder_Sum $T=19060 -16515 0 0 $X=29500 $Y=-36080
X15 Z<2> 23 22 20 21 24 19 15 52 GND 16 53 18 54 14 55 17 56 13 57
+ VDD
+ 6_FA_v3 $T=62150 -60875 0 0 $X=53915 $Y=-76150
X16 Z<3> 26 28 27 29 30 25 23 59 GND 22 60 20 61 21 62 24 63 19 64
+ VDD
+ 6_FA_v3 $T=86850 -60875 0 0 $X=78615 $Y=-76150
X17 Z<4> Z<5> Z<6> Z<7> Z<8> Z<9> Z<10> 26 66 GND 28 67 27 68 29 69 30 70 25 71
+ VDD
+ 6_FA_v3 $T=111575 -60875 0 0 $X=103340 $Y=-76150
X18 X<0> X<1> X<2> X<3> GND VDD Y<1> 7 8 Y<1> 9 10 ICV_3 $T=18540 -72855 0 90 $X=19065 $Y=-71875
X19 X<4> X<5> X<0> X<1> GND VDD Y<1> 11 12 Y<0> Z<0> 34 ICV_3 $T=18540 -60135 0 90 $X=19065 $Y=-59155
X20 X<2> X<3> X<4> X<5> GND VDD Y<0> 35 36 Y<0> 37 38 ICV_3 $T=18540 -47415 0 90 $X=19065 $Y=-46435
.ENDS
***************************************
