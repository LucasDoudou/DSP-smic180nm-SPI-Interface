* SPICE NETLIST
***************************************

.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_3 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_5 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_2 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_7 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_6 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_3 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_3 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_5 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_5 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_2 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_2 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_4 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_4 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_7 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_7 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_6 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_6 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=48
X0 1 6 5 2 8 9 7 Full_Adder_Sum $T=0 0 0 0 $X=10440 $Y=-19565
X1 3 11 10 4 8 9 12 Full_Adder_Sum $T=0 7690 0 0 $X=10440 $Y=-11875
.ENDS
***************************************
.SUBCKT 11FA_v3 COUT S<0> S<1> S<2> S<3> S<4> S<5> S<6> S<7> S<8> S<9> S<10> GND VDD B<6> A<6> B<7> A<7> B<10> A<10>
+ B<0> A<0> B<1> A<1> B<2> A<2> B<3> A<3> B<4> A<4> B<5> A<5> B<8> A<8> B<9> A<9>
** N=68 EP=36 IP=135 FDC=308
X0 36 GND VDD S<0> 1 27 ICV_1 $T=12585 -25495 0 0 $X=8470 $Y=-22410
X1 37 GND VDD S<1> 2 28 ICV_1 $T=12585 -17805 0 0 $X=8470 $Y=-14720
X2 38 GND VDD S<2> 3 29 ICV_1 $T=12585 -9930 0 0 $X=8470 $Y=-6845
X3 39 GND VDD S<3> 4 24 ICV_1 $T=12585 -2240 0 0 $X=8470 $Y=845
X4 40 GND VDD S<4> 5 30 ICV_1 $T=12585 5585 0 0 $X=8470 $Y=8670
X5 41 GND VDD S<5> 6 25 ICV_1 $T=12585 13275 0 0 $X=8470 $Y=16360
X6 42 GND VDD S<6> 7 31 ICV_1 $T=12585 20875 0 0 $X=8470 $Y=23960
X7 43 GND VDD S<7> 8 32 ICV_1 $T=12585 28405 0 0 $X=8470 $Y=31490
X8 44 GND VDD S<8> 9 33 ICV_1 $T=12585 36280 0 0 $X=8470 $Y=39365
X9 45 GND VDD S<9> 10 26 ICV_1 $T=12585 43970 0 0 $X=8470 $Y=47055
X10 46 GND VDD S<10> 11 COUT ICV_1 $T=12585 51795 0 0 $X=8470 $Y=54880
X11 25 A<6> B<6> 7 GND VDD 42 Full_Adder_Sum $T=-17040 43525 0 0 $X=-6600 $Y=23960
X12 31 A<7> B<7> 8 GND VDD 43 Full_Adder_Sum $T=-17040 51055 0 0 $X=-6600 $Y=31490
X13 26 A<10> B<10> 11 GND VDD 46 Full_Adder_Sum $T=-17040 74445 0 0 $X=-6600 $Y=54880
X14 GND 1 27 2 B<0> A<0> 36 GND VDD B<1> A<1> 37 ICV_2 $T=-17040 -2845 0 0 $X=-6600 $Y=-22410
X15 28 3 29 4 B<2> A<2> 38 GND VDD B<3> A<3> 39 ICV_2 $T=-17040 12720 0 0 $X=-6600 $Y=-6845
X16 24 5 30 6 B<4> A<4> 40 GND VDD B<5> A<5> 41 ICV_2 $T=-17040 28235 0 0 $X=-6600 $Y=8670
X17 32 9 33 10 B<8> A<8> 44 GND VDD B<9> A<9> 45 ICV_2 $T=-17040 58930 0 0 $X=-6600 $Y=39365
.ENDS
***************************************
