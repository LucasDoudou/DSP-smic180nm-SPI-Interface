* SPICE NETLIST
***************************************

.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT 4_Full_Adder_Type28 S<0> S<1> S<2> S<3> CO GND VDD B<0> A<0> B<1> A<1> B<2> A<2> B<3> A<3>
** N=26 EP=15 IP=60 FDC=112
X0 GND A<0> B<0> 1 GND VDD 15 Full_Adder_Sum $T=-8750 1760 0 0 $X=1690 $Y=-17805
X1 10 A<1> B<1> 2 GND VDD 16 Full_Adder_Sum $T=-8750 9450 0 0 $X=1690 $Y=-10115
X2 11 A<2> B<2> 3 GND VDD 17 Full_Adder_Sum $T=-8750 17325 0 0 $X=1690 $Y=-2240
X3 12 A<3> B<3> 4 GND VDD 18 Full_Adder_Sum $T=-8750 25015 0 0 $X=1690 $Y=5450
X4 15 GND VDD S<0> inv $T=20875 -20890 0 0 $X=16760 $Y=-17805
X5 16 GND VDD S<1> inv $T=20875 -13200 0 0 $X=16760 $Y=-10115
X6 17 GND VDD S<2> inv $T=20875 -5325 0 0 $X=16760 $Y=-2240
X7 18 GND VDD S<3> inv $T=20875 2365 0 0 $X=16760 $Y=5450
X8 1 GND VDD 10 inv $T=22375 -20890 0 0 $X=18260 $Y=-17805
X9 2 GND VDD 11 inv $T=22375 -13200 0 0 $X=18260 $Y=-10115
X10 3 GND VDD 12 inv $T=22375 -5325 0 0 $X=18260 $Y=-2240
X11 4 GND VDD CO inv $T=22375 2365 0 0 $X=18260 $Y=5450
.ENDS
***************************************
