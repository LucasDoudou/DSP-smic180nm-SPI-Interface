* SPICE NETLIST
***************************************

.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 5 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 12 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 8 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 11 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 5 VDD 5 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 10 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 8 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 9 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 12 VDD 12 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 11 GND 11 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
