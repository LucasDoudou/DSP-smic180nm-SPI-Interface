* SPICE NETLIST
***************************************

.SUBCKT inv_v2 VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=1410 $Y=-3310 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1410 $Y=-1870 $D=4
.ENDS
***************************************
