* SPICE NETLIST
***************************************

.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_3 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_5 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_2 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_7 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_6 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_3 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_3 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_5 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_5 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_2 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_2 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_4 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_4 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_7 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_7 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_6 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_6 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT And_Gate VIN_B VIN_A VDD GND VOUT
** N=7 EP=5 IP=0 FDC=6
M0 6 VIN_A 7 GND NM L=1.8e-07 W=2.2e-07 $X=1890 $Y=-4485 $D=0
M1 GND VIN_B 6 GND NM L=1.8e-07 W=2.2e-07 $X=2690 $Y=-4485 $D=0
M2 VOUT 7 GND GND NM L=1.8e-07 W=2.2e-07 $X=3490 $Y=-4485 $D=0
M3 7 VIN_A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1890 $Y=-2095 $D=4
M4 VDD VIN_B 7 VDD PM L=1.8e-07 W=4.4e-07 $X=2610 $Y=-2095 $D=4
M5 VOUT 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3330 $Y=-2095 $D=4
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=12
X0 1 3 5 4 6 And_Gate $T=0 0 0 0 $X=980 $Y=-5625
X1 2 3 5 4 7 And_Gate $T=3180 0 0 0 $X=4160 $Y=-5625
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=24
X0 1 2 5 6 7 8 9 ICV_2 $T=0 0 0 0 $X=980 $Y=-5625
X1 3 4 10 6 7 11 12 ICV_2 $T=6360 0 0 0 $X=7340 $Y=-5625
.ENDS
***************************************
.SUBCKT 5_6_Mul_draft2 X<0> X<1> X<2> X<3> X<4> X<5> Y<1> Y<0> Z<0> Z<1> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> GND VDD
** N=46 EP=18 IP=114 FDC=240
X0 41 GND VDD Z<1> 21 36 ICV_1 $T=46290 -55845 0 0 $X=42175 $Y=-52760
X1 42 GND VDD OUT<1> 22 37 ICV_1 $T=46290 -48155 0 0 $X=42175 $Y=-45070
X2 43 GND VDD OUT<2> 23 38 ICV_1 $T=46290 -40280 0 0 $X=42175 $Y=-37195
X3 44 GND VDD OUT<3> 24 35 ICV_1 $T=46290 -32590 0 0 $X=42175 $Y=-29505
X4 45 GND VDD OUT<4> 25 39 ICV_1 $T=46290 -24765 0 0 $X=42175 $Y=-21680
X5 46 GND VDD OUT<5> 26 OUT<6> ICV_1 $T=46290 -17075 0 0 $X=42175 $Y=-13990
X6 GND 16 7 21 GND VDD 41 Full_Adder_Sum $T=16665 -33195 0 0 $X=27105 $Y=-52760
X7 36 17 8 22 GND VDD 42 Full_Adder_Sum $T=16665 -25505 0 0 $X=27105 $Y=-45070
X8 37 18 9 23 GND VDD 43 Full_Adder_Sum $T=16665 -17630 0 0 $X=27105 $Y=-37195
X9 38 19 10 24 GND VDD 44 Full_Adder_Sum $T=16665 -9940 0 0 $X=27105 $Y=-29505
X10 35 20 11 25 GND VDD 45 Full_Adder_Sum $T=16665 -2115 0 0 $X=27105 $Y=-21680
X11 39 GND 12 26 GND VDD 46 Full_Adder_Sum $T=16665 5575 0 0 $X=27105 $Y=-13990
X12 X<0> X<1> X<2> X<3> Y<1> GND VDD 7 8 Y<1> 9 10 ICV_3 $T=16145 -50765 0 90 $X=16670 $Y=-49785
X13 X<4> X<5> X<0> X<1> Y<1> GND VDD 11 12 Y<0> Z<0> 16 ICV_3 $T=16145 -38045 0 90 $X=16670 $Y=-37065
X14 X<2> X<3> X<4> X<5> Y<0> GND VDD 17 18 Y<0> 19 20 ICV_3 $T=16145 -25325 0 90 $X=16670 $Y=-24345
.ENDS
***************************************
