* SPICE NETLIST
***************************************

.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_3 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_5 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_2 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_7 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_6 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_3 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_3 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_5 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_5 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_2 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_2 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_4 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_4 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_7 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_7 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_6 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_6 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=48
X0 1 2 3 4 10 11 9 Full_Adder_Sum $T=0 0 0 0 $X=10440 $Y=-19565
X1 5 6 7 8 10 11 12 Full_Adder_Sum $T=0 7690 0 0 $X=10440 $Y=-11875
.ENDS
***************************************
.SUBCKT 11FA_v4 B<0> B<1> B<2> B<3> B<4> B<5> A<0> A<1> A<2> A<3> A<4> A<5> S<1> S<2> S<3> S<4> S<5> S<0> B<9> A<7>
+ A<8> B<10> A<6> B<6> A<9> A<10> B<8> B<7> S<6> S<7> S<8> S<9> S<10> COUT GND VDD
** N=68 EP=36 IP=133 FDC=308
X0 58 GND VDD S<0> 36 43 ICV_1 $T=26880 -61070 0 0 $X=22765 $Y=-57985
X1 59 GND VDD S<1> 37 44 ICV_1 $T=26880 -53380 0 0 $X=22765 $Y=-50295
X2 60 GND VDD S<2> 38 45 ICV_1 $T=26880 -45505 0 0 $X=22765 $Y=-42420
X3 61 GND VDD S<3> 39 42 ICV_1 $T=26880 -37815 0 0 $X=22765 $Y=-34730
X4 62 GND VDD S<4> 40 46 ICV_1 $T=26880 -29990 0 0 $X=22765 $Y=-26905
X5 63 GND VDD S<5> 41 18 ICV_1 $T=26880 -22300 0 0 $X=22765 $Y=-19215
X6 64 GND VDD S<6> 47 52 ICV_1 $T=47180 -53190 0 0 $X=43065 $Y=-50105
X7 65 GND VDD S<7> 48 53 ICV_1 $T=47180 -45500 0 0 $X=43065 $Y=-42415
X8 66 GND VDD S<8> 49 54 ICV_1 $T=47180 -37625 0 0 $X=43065 $Y=-34540
X9 67 GND VDD S<9> 50 55 ICV_1 $T=47180 -29935 0 0 $X=43065 $Y=-26850
X10 68 GND VDD S<10> 51 COUT ICV_1 $T=47180 -22300 0 0 $X=43065 $Y=-19215
X11 55 A<10> B<10> 51 GND VDD 68 Full_Adder_Sum $T=17555 350 0 0 $X=27995 $Y=-19215
X12 GND A<0> B<0> 36 43 A<1> B<1> 37 58 GND VDD 59 ICV_2 $T=-2745 -38420 0 0 $X=7695 $Y=-57985
X13 44 A<2> B<2> 38 45 A<3> B<3> 39 60 GND VDD 61 ICV_2 $T=-2745 -22855 0 0 $X=7695 $Y=-42420
X14 42 A<4> B<4> 40 46 A<5> B<5> 41 62 GND VDD 63 ICV_2 $T=-2745 -7340 0 0 $X=7695 $Y=-26905
X15 18 A<6> B<6> 47 52 A<7> B<7> 48 64 GND VDD 65 ICV_2 $T=17555 -30540 0 0 $X=27995 $Y=-50105
X16 53 A<8> B<8> 49 54 A<9> B<9> 50 66 GND VDD 67 ICV_2 $T=17555 -14975 0 0 $X=27995 $Y=-34540
.ENDS
***************************************
