* SPICE NETLIST
***************************************

.SUBCKT And_Gate VIN_B VIN_A VDD GND VOUT
** N=7 EP=5 IP=0 FDC=6
M0 6 VIN_A 7 GND NM L=1.8e-07 W=2.2e-07 $X=1890 $Y=-4485 $D=0
M1 GND VIN_B 6 GND NM L=1.8e-07 W=2.2e-07 $X=2690 $Y=-4485 $D=0
M2 VOUT 7 GND GND NM L=1.8e-07 W=2.2e-07 $X=3490 $Y=-4485 $D=0
M3 7 VIN_A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1890 $Y=-2095 $D=4
M4 VDD VIN_B 7 VDD PM L=1.8e-07 W=4.4e-07 $X=2610 $Y=-2095 $D=4
M5 VOUT 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3330 $Y=-2095 $D=4
.ENDS
***************************************
.SUBCKT 6_AND_test Y<0> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND Z<0> A<0> A<1> A<2> A<3> A<4>
** N=15 EP=15 IP=30 FDC=36
X0 X<0> Y<0> VDD GND Z<0> And_Gate $T=2375 -2105 0 0 $X=3355 $Y=-7730
X1 X<1> Y<0> VDD GND A<0> And_Gate $T=5555 -2105 0 0 $X=6535 $Y=-7730
X2 X<2> Y<0> VDD GND A<1> And_Gate $T=8735 -2105 0 0 $X=9715 $Y=-7730
X3 X<3> Y<0> VDD GND A<2> And_Gate $T=11915 -2105 0 0 $X=12895 $Y=-7730
X4 X<4> Y<0> VDD GND A<3> And_Gate $T=15095 -2105 0 0 $X=16075 $Y=-7730
X5 X<5> Y<0> VDD GND A<4> And_Gate $T=18275 -2105 0 0 $X=19255 $Y=-7730
.ENDS
***************************************
.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT 6_FA_v3 S<0> S<1> S<2> S<3> S<4> S<5> S<6> A<0> B<0> GND A<1> B<1> A<2> B<2> A<3> B<3> A<4> B<4> A<5> B<5>
+ VDD
** N=38 EP=21 IP=78 FDC=168
X0 33 GND VDD S<0> 22 29 ICV_1 $T=11635 -18360 0 0 $X=7520 $Y=-15275
X1 34 GND VDD S<1> 23 30 ICV_1 $T=11635 -10670 0 0 $X=7520 $Y=-7585
X2 35 GND VDD S<2> 24 31 ICV_1 $T=11635 -2795 0 0 $X=7520 $Y=290
X3 36 GND VDD S<3> 25 28 ICV_1 $T=11635 4895 0 0 $X=7520 $Y=7980
X4 37 GND VDD S<4> 26 32 ICV_1 $T=11635 12720 0 0 $X=7520 $Y=15805
X5 38 GND VDD S<5> 27 S<6> ICV_1 $T=11635 20410 0 0 $X=7520 $Y=23495
X6 GND A<0> B<0> 22 GND VDD 33 Full_Adder_Sum $T=-17990 4290 0 0 $X=-7550 $Y=-15275
X7 29 A<1> B<1> 23 GND VDD 34 Full_Adder_Sum $T=-17990 11980 0 0 $X=-7550 $Y=-7585
X8 30 A<2> B<2> 24 GND VDD 35 Full_Adder_Sum $T=-17990 19855 0 0 $X=-7550 $Y=290
X9 31 A<3> B<3> 25 GND VDD 36 Full_Adder_Sum $T=-17990 27545 0 0 $X=-7550 $Y=7980
X10 28 A<4> B<4> 26 GND VDD 37 Full_Adder_Sum $T=-17990 35370 0 0 $X=-7550 $Y=15805
X11 32 A<5> B<5> 27 GND VDD 38 Full_Adder_Sum $T=-17990 43060 0 0 $X=-7550 $Y=23495
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=12
X0 1 3 4 5 6 And_Gate $T=0 0 0 0 $X=980 $Y=-5625
X1 2 3 4 5 7 And_Gate $T=3180 0 0 0 $X=4160 $Y=-5625
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=24
X0 1 2 7 6 5 8 9 ICV_2 $T=0 0 0 0 $X=980 $Y=-5625
X1 3 4 10 6 5 11 12 ICV_2 $T=6360 0 0 0 $X=7340 $Y=-5625
.ENDS
***************************************
.SUBCKT 5_6_Mul_final_test1 X<0> X<1> X<2> X<3> X<4> X<5> Y<1> Y<0> Z<0> Z<1> GND Y<2> Y<3> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> VDD
+ Z<2> Z<3>
** N=74 EP=22 IP=186 FDC=648
X0 Y<2> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 47 48 49 50 51 52 6_AND_test $T=52435 -7615 0 0 $X=55595 $Y=-15345
X1 Y<3> X<0> X<1> X<2> X<3> X<4> X<5> VDD GND 54 55 56 57 58 59 6_AND_test $T=77135 -7615 0 0 $X=80295 $Y=-15345
X2 67 GND VDD Z<1> 33 42 ICV_1 $T=50010 -63130 0 0 $X=45895 $Y=-60045
X3 68 GND VDD 15 34 43 ICV_1 $T=50010 -55440 0 0 $X=45895 $Y=-52355
X4 69 GND VDD 16 35 44 ICV_1 $T=50010 -47565 0 0 $X=45895 $Y=-44480
X5 70 GND VDD 18 36 41 ICV_1 $T=50010 -39875 0 0 $X=45895 $Y=-36790
X6 71 GND VDD 14 37 45 ICV_1 $T=50010 -32050 0 0 $X=45895 $Y=-28965
X7 72 GND VDD 17 38 13 ICV_1 $T=50010 -24360 0 0 $X=45895 $Y=-21275
X8 GND 28 7 33 GND VDD 67 Full_Adder_Sum $T=20385 -40480 0 0 $X=30825 $Y=-60045
X9 42 29 8 34 GND VDD 68 Full_Adder_Sum $T=20385 -32790 0 0 $X=30825 $Y=-52355
X10 43 30 9 35 GND VDD 69 Full_Adder_Sum $T=20385 -24915 0 0 $X=30825 $Y=-44480
X11 44 31 10 36 GND VDD 70 Full_Adder_Sum $T=20385 -17225 0 0 $X=30825 $Y=-36790
X12 41 32 11 37 GND VDD 71 Full_Adder_Sum $T=20385 -9400 0 0 $X=30825 $Y=-28965
X13 45 GND 12 38 GND VDD 72 Full_Adder_Sum $T=20385 -1710 0 0 $X=30825 $Y=-21275
X14 Z<2> 23 22 20 21 24 19 15 47 GND 16 48 18 49 14 50 17 51 13 52
+ VDD
+ 6_FA_v3 $T=63475 -46070 0 0 $X=55240 $Y=-61345
X15 Z<3> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> 23 54 GND 22 55 20 56 21 57 24 58 19 59
+ VDD
+ 6_FA_v3 $T=88175 -46070 0 0 $X=79940 $Y=-61345
X16 X<0> X<1> X<2> X<3> GND VDD Y<1> 7 8 Y<1> 9 10 ICV_3 $T=19865 -58050 0 90 $X=20390 $Y=-57070
X17 X<4> X<5> X<0> X<1> GND VDD Y<1> 11 12 Y<0> Z<0> 28 ICV_3 $T=19865 -45330 0 90 $X=20390 $Y=-44350
X18 X<2> X<3> X<4> X<5> GND VDD Y<0> 29 30 Y<0> 31 32 ICV_3 $T=19865 -32610 0 90 $X=20390 $Y=-31630
.ENDS
***************************************
