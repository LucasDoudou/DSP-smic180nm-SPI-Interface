* SPICE NETLIST
***************************************

.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=48
X0 1 2 3 4 10 11 9 Full_Adder_Sum $T=0 0 0 0 $X=10440 $Y=-19565
X1 5 6 7 8 10 11 12 Full_Adder_Sum $T=0 7690 0 0 $X=10440 $Y=-11875
.ENDS
***************************************
.SUBCKT 11FA_v1 B<9> A<7> A<8> B<10> A<6> B<6> A<9> A<10> B<8> B<7> S<5> S<1> S<2> S<3> S<4> S<0> S<6> S<7> S<8> S<9>
+ S<10> COUT GND A<1> B<1> A<0> B<0> A<3> B<3> A<2> B<2> A<5> B<5> A<4> B<4> VDD
** N=68 EP=36 IP=133 FDC=308
X0 58 GND VDD S<0> 11 20 ICV_1 $T=11565 -26110 0 0 $X=7450 $Y=-23025
X1 59 GND VDD S<1> 12 21 ICV_1 $T=11565 -18420 0 0 $X=7450 $Y=-15335
X2 60 GND VDD S<2> 13 22 ICV_1 $T=11565 -10545 0 0 $X=7450 $Y=-7460
X3 61 GND VDD S<3> 14 19 ICV_1 $T=11565 -2855 0 0 $X=7450 $Y=230
X4 62 GND VDD S<4> 15 23 ICV_1 $T=11565 4970 0 0 $X=7450 $Y=8055
X5 63 GND VDD S<5> 16 18 ICV_1 $T=11565 12660 0 0 $X=7450 $Y=15745
X6 64 GND VDD S<6> 29 40 ICV_1 $T=35330 -18230 0 0 $X=31215 $Y=-15145
X7 65 GND VDD S<7> 30 41 ICV_1 $T=35330 -10540 0 0 $X=31215 $Y=-7455
X8 66 GND VDD S<8> 31 42 ICV_1 $T=35330 -2665 0 0 $X=31215 $Y=420
X9 67 GND VDD S<9> 32 43 ICV_1 $T=35330 5025 0 0 $X=31215 $Y=8110
X10 68 GND VDD S<10> 33 COUT ICV_1 $T=35330 12660 0 0 $X=31215 $Y=15745
X11 43 A<10> B<10> 33 GND VDD 68 Full_Adder_Sum $T=5705 35310 0 0 $X=16145 $Y=15745
X12 GND A<0> B<0> 11 20 A<1> B<1> 12 58 GND VDD 59 ICV_2 $T=-18060 -3460 0 0 $X=-7620 $Y=-23025
X13 21 A<2> B<2> 13 22 A<3> B<3> 14 60 GND VDD 61 ICV_2 $T=-18060 12105 0 0 $X=-7620 $Y=-7460
X14 19 A<4> B<4> 15 23 A<5> B<5> 16 62 GND VDD 63 ICV_2 $T=-18060 27620 0 0 $X=-7620 $Y=8055
X15 18 A<6> B<6> 29 40 A<7> B<7> 30 64 GND VDD 65 ICV_2 $T=5705 4420 0 0 $X=16145 $Y=-15145
X16 41 A<8> B<8> 31 42 A<9> B<9> 32 66 GND VDD 67 ICV_2 $T=5705 19985 0 0 $X=16145 $Y=420
.ENDS
***************************************
