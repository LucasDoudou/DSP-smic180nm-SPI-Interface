* SPICE NETLIST
***************************************

.SUBCKT inv VI GND VDD VO
** N=4 EP=4 IP=0 FDC=2
M0 VO VI GND GND NM L=1.8e-07 W=2.2e-07 $X=-3205 $Y=4225 $D=0
M1 VO VI VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-3205 $Y=5665 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 4 inv $T=0 0 0 0 $X=-4115 $Y=3085
X1 5 2 3 6 inv $T=1500 0 0 0 $X=-2615 $Y=3085
.ENDS
***************************************
.SUBCKT And_Gate VIN_B VIN_A VDD GND VOUT
** N=7 EP=5 IP=0 FDC=6
M0 6 VIN_A 7 GND NM L=1.8e-07 W=2.2e-07 $X=1890 $Y=-4485 $D=0
M1 GND VIN_B 6 GND NM L=1.8e-07 W=2.2e-07 $X=2690 $Y=-4485 $D=0
M2 VOUT 7 GND GND NM L=1.8e-07 W=2.2e-07 $X=3490 $Y=-4485 $D=0
M3 7 VIN_A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=1890 $Y=-2095 $D=4
M4 VDD VIN_B 7 VDD PM L=1.8e-07 W=4.4e-07 $X=2610 $Y=-2095 $D=4
M5 VOUT 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3330 $Y=-2095 $D=4
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=12
X0 1 3 5 4 6 And_Gate $T=0 0 0 0 $X=980 $Y=-5625
X1 2 3 5 4 7 And_Gate $T=3180 0 0 0 $X=4160 $Y=-5625
.ENDS
***************************************
.SUBCKT p18_1 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_3 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_0 1 2 3 4 5 6
** N=7 EP=6 IP=0 FDC=2
M0 3 5 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 6 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_2 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 1 5 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_5 1 2 3 4 5 6 7 8
** N=9 EP=8 IP=0 FDC=3
M0 3 6 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
M1 4 7 3 1 PM L=1.8e-07 W=8.8e-07 $X=720 $Y=0 $D=4
M2 5 8 4 1 PM L=1.8e-07 W=8.8e-07 $X=1440 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=0 FDC=3
M0 3 6 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
M1 4 7 3 1 NM L=1.8e-07 W=4.4e-07 $X=720 $Y=0 $D=0
M2 5 8 4 1 NM L=1.8e-07 W=4.4e-07 $X=1440 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Full_Adder_Sum CI A B CO_ GND VDD S_
** N=17 EP=7 IP=76 FDC=24
X0 VDD CO_ 8 CI p18_1 $T=11350 -14410 0 0 $X=10440 $Y=-14840
X1 VDD S_ 13 CO_ p18_1 $T=17285 -14410 0 0 $X=16375 $Y=-14840
X2 GND CO_ 9 CI n18_3 $T=11350 -18435 0 0 $X=10690 $Y=-19565
X3 GND S_ 12 CO_ n18_3 $T=17285 -18435 0 0 $X=16625 $Y=-19565
X4 VDD 8 VDD 8 B A p18_0 $T=12845 -14410 0 0 $X=11935 $Y=-14840
X5 VDD CO_ 11 VDD B A p18_0 $T=15065 -14410 0 0 $X=14155 $Y=-14840
X6 GND GND 9 B A n18_2 $T=12845 -18435 0 0 $X=12185 $Y=-19565
X7 GND CO_ 10 B A n18_2 $T=15065 -18435 0 0 $X=14405 $Y=-19565
X8 VDD VDD 13 VDD 13 CI A B p18_5 $T=18785 -14410 0 0 $X=17875 $Y=-14840
X9 VDD S_ 14 17 VDD CI A B p18_5 $T=21725 -14410 0 0 $X=20815 $Y=-14840
X10 GND GND 12 GND 12 CI A B n18_4 $T=18785 -18435 0 0 $X=18125 $Y=-19565
X11 GND S_ 15 16 GND CI A B n18_4 $T=21725 -18435 0 0 $X=21065 $Y=-19565
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=48
X0 3 1 2 4 9 10 11 Full_Adder_Sum $T=0 0 0 0 $X=10440 $Y=-19565
X1 7 5 6 8 9 10 12 Full_Adder_Sum $T=0 7690 0 0 $X=10440 $Y=-11875
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=24
X0 1 2 5 6 7 8 9 ICV_2 $T=0 0 0 0 $X=980 $Y=-5625
X1 3 4 10 6 7 11 12 ICV_2 $T=6360 0 0 0 $X=7340 $Y=-5625
.ENDS
***************************************
.SUBCKT 5_6_Mul_draft1 X<0> X<1> X<2> X<3> X<4> X<5> Y<1> Y<0> Z<0> Z<1> GND Y<2> Z<2> OUT3<1> OUT3<2> OUT3<3> OUT3<4> OUT3<5> OUT3<6> VDD
** N=77 EP=20 IP=201 FDC=444
X0 66 GND VDD Z<1> 27 36 ICV_1 $T=50010 -63130 0 0 $X=45895 $Y=-60045
X1 67 GND VDD 15 28 37 ICV_1 $T=50010 -55440 0 0 $X=45895 $Y=-52355
X2 68 GND VDD 16 29 38 ICV_1 $T=50010 -47565 0 0 $X=45895 $Y=-44480
X3 69 GND VDD 18 30 35 ICV_1 $T=50010 -39875 0 0 $X=45895 $Y=-36790
X4 70 GND VDD 14 31 39 ICV_1 $T=50010 -32050 0 0 $X=45895 $Y=-28965
X5 71 GND VDD 17 32 13 ICV_1 $T=50010 -24360 0 0 $X=45895 $Y=-21275
X6 72 GND VDD Z<2> 46 60 ICV_1 $T=75110 -64430 0 0 $X=70995 $Y=-61345
X7 73 GND VDD OUT3<1> 47 61 ICV_1 $T=75110 -56740 0 0 $X=70995 $Y=-53655
X8 74 GND VDD OUT3<2> 48 62 ICV_1 $T=75110 -48865 0 0 $X=70995 $Y=-45780
X9 75 GND VDD OUT3<3> 49 59 ICV_1 $T=75110 -41175 0 0 $X=70995 $Y=-38090
X10 76 GND VDD OUT3<4> 50 63 ICV_1 $T=75110 -33350 0 0 $X=70995 $Y=-30265
X11 77 GND VDD OUT3<5> 51 OUT3<6> ICV_1 $T=75110 -25660 0 0 $X=70995 $Y=-22575
X12 X<0> X<1> Y<2> GND VDD 40 41 ICV_2 $T=54810 -9720 0 0 $X=55790 $Y=-15345
X13 X<2> X<3> Y<2> GND VDD 42 43 ICV_2 $T=61170 -9720 0 0 $X=62150 $Y=-15345
X14 X<4> X<5> Y<2> GND VDD 44 64 ICV_2 $T=67530 -9720 0 0 $X=68510 $Y=-15345
X15 22 7 GND 27 23 8 36 28 GND VDD 66 67 ICV_3 $T=20385 -40480 0 0 $X=30825 $Y=-60045
X16 24 9 37 29 25 10 38 30 GND VDD 68 69 ICV_3 $T=20385 -24915 0 0 $X=30825 $Y=-44480
X17 26 11 35 31 GND 12 39 32 GND VDD 70 71 ICV_3 $T=20385 -9400 0 0 $X=30825 $Y=-28965
X18 15 40 GND 46 16 41 60 47 GND VDD 72 73 ICV_3 $T=45485 -41780 0 0 $X=55925 $Y=-61345
X19 18 42 61 48 14 43 62 49 GND VDD 74 75 ICV_3 $T=45485 -26215 0 0 $X=55925 $Y=-45780
X20 17 44 59 50 13 64 63 51 GND VDD 76 77 ICV_3 $T=45485 -10700 0 0 $X=55925 $Y=-30265
X21 X<0> X<1> X<2> X<3> Y<1> GND VDD 7 8 Y<1> 9 10 ICV_4 $T=19865 -58050 0 90 $X=20390 $Y=-57070
X22 X<4> X<5> X<0> X<1> Y<1> GND VDD 11 12 Y<0> Z<0> 22 ICV_4 $T=19865 -45330 0 90 $X=20390 $Y=-44350
X23 X<2> X<3> X<4> X<5> Y<0> GND VDD 23 24 Y<0> 25 26 ICV_4 $T=19865 -32610 0 90 $X=20390 $Y=-31630
.ENDS
***************************************
